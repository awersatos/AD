* SPICE MODEL LMV711
* BEGIN MODEL
.SUBCKT LMV711  8 42 1 24 25 30
* PINOUT ORDER +IN -IN V+ V- OUT SD
*               8   42  1 24  25 30
C5 0 29 10.0E-12
E4 21 15 8 15 0.5
R1 1 11 4.8E3
C6 42 0 10.0E-12
R2 1 12 4.8E3
R3 9 24 4.8E3
R4 10 24 4.8E3
G1 15 16 11 12 145.0E-6
G2 15 16 9 10 145.0E-6
R5 1 17 10.0E6
R6 17 24 10.0E6
E1 15 0 17 0 1.0
R7 16 15 50.7E6
V3 1 20 1.37
V4 18 24 1.37
I2 22 23 10.0E-6
I3 26 13 10.0E-6
C1 16 25 2.5E-12
E2 31 24 16 15 1.0
E3 1 47 15 16 1.0
R11 36 24 15.5
R12 1 35 20.0
R13 32 35 1.0E3
E5 28 21 42 15 0.5
R9 28 27 1.0E6
C2 28 27 0.75E-12
R10 27 15 10.0E3
E6 8 29 27 15 1.0E-3
C7 29 42 4.0E-12
C8 11 12 1.5E-12
R14 33 36 1.0E3
C9 9 10 1.5E-12
D9 13 26 D1M
E7 23 36 48 22 100.0
VIQ 69 0 8.0
G6 1 24 68 24 100.0E-6
RIQ 68 69 100.0E6
R16 22 36 1.0E3
E8 26 35 19 13 100.0
R17 35 13 1.0E3
R22 30 40 400.0
G3 1 3 6 24 1.0E-6
V8 43 24 21.65
R15 43 6 1.0E6
C3 40 24 10.0E-12
R18 47 19 1.0E3
R19 31 48 1.0E3
G4 38 13 4 24 1.0E-6
V14 50 24 132.0
R20 50 4 1.0E6
G5 22 37 51 24 1.0E-6
V15 54 24 132.0
R21 54 51 1.0E6
V16 41 24 1.3
V17 1 7 1.37
V18 14 42 300.0E-6
V19 42 44 200.0E-6
D1 16 20 D1M
D2 18 16 D1M
D3 2 1 D1M
D4 8 1 D1M
D5 24 8 D1M
D6 24 44 D1M
D7 14 1 D1M
D8 23 22 D1M
Q1 16 32 1 NBJT
Q2 16 33 24 PBJT
MIQ 68 39 24 24 M10M L=6U W=6U
M1 34 53 1 1 M1M L=6U W=100U
M5 11 29 5 24 M2M L=6U W=25U
M6 12 14 5 24 M2M L=6U W=25U
M7 9 29 2 2 M1M L=6U W=25U
M8 10 42 2 2 M1M L=6U W=25U
M9 25 38 35 35 M9M L=1.5U W=500U
M10 25 37 36 36 NOX L=1.5U W=500U
M13 37 37 22 22 NOX L=1.5U W=500U
M14 38 38 13 13 M9M L=1.5U W=500U
M15 37 39 24 24 M3M L=6U W=6U
M16 38 40 1 1 M4M L=6U W=6U
M17 39 40 1 1 M4M L=6U W=0.6U
M18 39 40 24 24 M3M L=6U W=0.6U
M19 6 39 24 24 M3M L=6U W=6U
M20 25 39 24 24 M7M L=1.5U W=500U
M21 19 40 1 1 M4M L=6U W=6U
M22 48 39 24 24 M3M L=6U W=6U
M23 4 39 24 24 M3M L=6U W=6U
M24 51 39 24 24 M3M L=6U W=6U
M25 2 7 34 1 M1M L=6U W=100U
M26 3 3 24 24 M2M L=6U W=100U
M27 53 41 5 5 M2M L=6U W=100U
M28 5 3 24 24 M2M L=6U W=100U
M30 53 53 1 1 M1M L=6U W=100U
.MODEL D1M D CJO=0.1E-12
.MODEL NBJT PNP
.MODEL PBJT NPN
.MODEL M9M PMOS CBD=0.2E-12 CBS=0.2E-12 CGBO=50E-9
+ CGDO=50E-12 CGSO=50E-12 KP=200U LAMBDA=0.07
+ RD=1.0 RS=1.0 VTO=-0.75
.MODEL NOX NMOS CBD=0.2E-12 CBS=0.2E-12 CGBO=50E-9
+ CGDO=50e-12 CGSO=50e-12 KP=200u LAMBDA=0.07
+ RD=1.0 RS=1.0 VTO=0.75
.MODEL M1M PMOS KP=200U RD=1.0 RS=1.0 VTO=-0.75
.MODEL M2M NMOS KP=200U RD=1.0 RS=1.0 VTO=0.75
.MODEL M3M NMOS CBD=0.2E-12 CBS=0.2E-12 CGBO=10E-9
+ CGDO=5E-9 CGSO=5E-9 KP=200U RD=1.0 RS=1.0 VTO=0.75
.MODEL M4M PMOS CBD=0.2E-12 CBS=0.2E-12 CGBO=10E-9
+ CGDO=5E-9 CGSO=5E-9 KP=200U RD=1.0 RS=1.0 VTO=-0.75
.MODEL M10M NMOS CBD=0.2E-12 CBS=0.2E-12 CGBO=10E-9
+ CGDO=5E-9 CGSO=5E-9 KP=200U IS=1E-16 RS=1.0 VTO=0.75
.MODEL M7M NMOS CBD=0.2E-12 CBS=0.2E-12 CGBO=50E-9
+ CGDO=50E-12 CGSO=50E-12 KP=200U
+ RD=1.0 RS=1.0 VTO=1.75
.ENDS

