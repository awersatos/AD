*Default SCR
*SCR - pin order: A G K
.SUBCKT SCR  1 2 3
Q1 2 4 1 QPSCR AREA=.67 OFF
Q2 4 2 3 QNSCR AREA=.67
Q3 5 4 1 QPSCR AREA=.33 OFF
Q4 4 5 3 QNSCR AREA=.33
RBN 2 5 40
.MODEL QNSCR NPN(TF=400NS TR=1.6US CJC=75PF CJE=175PF XTB=2.5
+ IS=1E-14 ISE=3E-9 NE=2 BF=100 BR=25 ISC=3E-9 NC=2)
.MODEL QPSCR PNP(TF=90NS TR=180NS CJC=75PF CJE=80PF XTB=2.5 
+ IS=1E-14 ISE=3E-9 NE=2 BF=50 BR=25 ISC=3E-9 NC=2 RE=.03)
.ENDS SCR