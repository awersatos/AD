*IRF1010 MCE 4-2-96
*55V  75A .014 ohm HEXFET pkg:TO-220 2,1,3
.SUBCKT IRF1010  10 20 40 40
M1   1  2  3  3  DMOS L=1U W=1U
RD  10  1  5.65M
RS  30  3  1.35M
RG  20  2  12.1
CGS  2  3  2.15N
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  4.49N
R1  13  0  1
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.5N
.MODEL DMOS NMOS (LEVEL=3 THETA=60M VMAX=114K ETA=2M VTO=3 KP=19.4)
.MODEL DCGD D (CJO=4.49N VJ=.6 M=.68)
.MODEL DSUB D (IS=311N N=1.5 RS=8.67M BV=55 CJO=4.08N VJ=.8 M=.42 TT=100N)
.MODEL DLIM D (IS=100U)
.ENDS IRF1010

