-- "$Header: 42mx.vhd@@/main/4 $"
-- Actel Vital 95 library
library IEEE;
use IEEE.STD_LOGIC_1164.all;

library IEEE;
use IEEE.VITAL_Timing.all;

package COMPONENTS is

constant DefaultTimingChecksOn : Boolean := True;
constant DefaultXGenerationOn : Boolean := False;
constant DefaultXon : Boolean := False;
constant DefaultMsgOn : Boolean := True;

component AND2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND3C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND4B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND4C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND4D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AND5B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO10
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO11
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO1D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO1E
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO2C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO2D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO2E
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO3C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO5A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO6
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO6A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO7
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO8
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AO9
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI1D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AOI4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AX1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AX1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AX1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component AX1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component BBDLHS
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_GOUT_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_GIN_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_GOUT_noedge_negedge           :	VitalDelayType := 0.000 ns;
      tsetup_D_GOUT_noedge_negedge          :	VitalDelayType := 0.000 ns;
      thold_PAD_GIN_noedge_posedge          :	VitalDelayType := 0.000 ns;
      tsetup_PAD_GIN_noedge_posedge         :	VitalDelayType := 0.000 ns;
      tperiod_GIN_posedge            :	VitalDelayType := 0.000 ns;
      tperiod_GOUT_negedge           :	VitalDelayType := 0.000 ns;
      tpw_GIN_negedge                :	VitalDelayType := 0.000 ns;
      tpw_GOUT_posedge               :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_GIN                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_GOUT                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      GIN                            :	in    STD_ULOGIC;
      GOUT                           :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component BBHS
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component BIBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component BUFA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component BUFD
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component BUFF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CLKBIBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CLKBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CLKINT
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CM7
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S11_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S10_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CM8
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S11_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S10_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S01_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S00_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S00                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S01                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S00                            :	in    STD_ULOGIC;
      S01                            :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CS1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CS2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CY2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      A1                             :	in    STD_ULOGIC;
      B0                             :	in    STD_ULOGIC;
      B1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component CY2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      A1                             :	in    STD_ULOGIC;
      B0                             :	in    STD_ULOGIC;
      B1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component DF1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DF1_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DF1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DF1A_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DF1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DF1B_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DF1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DF1C_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFC1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1A_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1B_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1D_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFC1E
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFC1G
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFE
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE1B_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE1C_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE3C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFE3D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFEA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFEA_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFM1B_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFM1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFM1C_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFM3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM3E
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM4C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFM4D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFM6A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S1_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S1_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM6B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S1_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S1_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM7A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S10_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S10_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_S11_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S11_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFM7B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S10_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S10_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_S11_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S11_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFMA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFMA_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFMB
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFME1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1A_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1B_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFP1D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1D_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFP1E
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFP1F
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFP1G
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DFPC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFPC_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFPCA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DFPCA_CC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DL1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DL1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DL1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DL1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DL2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DL2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DL2C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DL2D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DLC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLC1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLC1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLC1F
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DLC1G
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DLCA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLE
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_E_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLE1D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DLE2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_CLR_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_CLR_E_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLE2C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_CLR_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_CLR_E_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLE3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_PRE_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_PRE_E_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLE3C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_PRE_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_PRE_E_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLEA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLEB
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_E_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLEC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_A_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_B                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_A_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_B                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S1_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S1_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S1_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S1_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S10_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S11_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S10_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S10_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S11_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S11_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLM4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S10_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S11_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S10_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S10_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S11_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S11_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLMA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLME1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_A_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_A_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_B_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_B_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_S_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLP1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLP1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLP1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLP1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component DLP1D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DLP1E
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component DXAND7
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_F_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_F                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      F                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component DXAX7
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_H_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_F_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_F                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_H                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      F                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      H                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component DXNAND7
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_F_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_F                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      F                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component FA1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CI_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CI_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CI                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CI                             :	in    STD_ULOGIC;
      S                              :	out   STD_ULOGIC;
      CO                             :	out   STD_ULOGIC);
end component; 

component FA1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CI_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CI_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CI                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CI                             :	in    STD_ULOGIC;
      S                              :	out   STD_ULOGIC;
      CO                             :	out   STD_ULOGIC);
end component; 

component FA2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CI_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CI_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CI                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      A1                             :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CI                             :	in    STD_ULOGIC;
      S                              :	out   STD_ULOGIC;
      CO                             :	out   STD_ULOGIC);
end component; 

component GAND2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component GMX4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component GNAND2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component GND
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True);

   port(
      Y                              :	out   STD_ULOGIC := '0');
end component; 

component GNOR2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component GOR2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component GXOR2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component HA1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
end component; 

component HA1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
end component; 

component HA1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
end component; 

component HA1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
end component; 

component IBDL
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_PAD_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_PAD_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component INBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component INV
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component INVA
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component INVD
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component IR
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_PAD_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_PAD_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component IRI
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_PAD_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_PAD_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
end component; 

component JKF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component JKF1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component JKF2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component JKF2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component JKF2C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component JKF2D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component MAJ3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component MX2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component MX2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component MX2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component MX2C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component MX4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component MXC1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component MXT
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0B_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0A_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0A                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0B                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0A                            :	in    STD_ULOGIC;
      S0B                            :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND3C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND4B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND4C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND4D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NAND5C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR3C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR4B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR4C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR4D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component NOR5C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA1C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OA5
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OAI1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OAI2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OAI3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OAI3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OBDLHS
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component OBHS
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component OR2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR2A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR2B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR3
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR3A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR3B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR3C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR4
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR4A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR4B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR4C
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR4D
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component OR5B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component ORH
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component ORIH
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component ORITH
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component ORTH
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component OUTBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component QCLKBUF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component QCLKINT
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component RAM4FA
  GENERIC (
        tipd_RDAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RDAD5_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD5_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD5_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD5_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_WRAD5_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  
end component; 

component RAM4FF
  GENERIC (
        tipd_RDAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD5_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  
end component; 

component RAM4FR
  GENERIC (
        tipd_RDAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD5_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  
end component; 

component RAM4RA
  GENERIC (
        tipd_RDAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RDAD5_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD5_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD5_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD5_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_WRAD5_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  
end component; 

component RAM4RF
  GENERIC (
        tipd_RDAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD5_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  
end component; 

component RAM4RR
  GENERIC (
        tipd_RDAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD5_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  
end component; 

component RAM8FA
  GENERIC (
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD7      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD6      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD5      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD4      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RDAD4_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_WRAD4_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC;
        RD6    : OUT STD_ULOGIC;
        RD5    : OUT STD_ULOGIC;
        RD4    : OUT STD_ULOGIC;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  
end component; 

component RAM8FF
  GENERIC (
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD7      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD6      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD5      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD4      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD4_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC;
        RD6    : OUT STD_ULOGIC;
        RD5    : OUT STD_ULOGIC;
        RD4    : OUT STD_ULOGIC;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  
end component; 

component RAM8FR
  GENERIC (
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD7      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD6      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD5      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD4      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD4_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC;
        RD6    : OUT STD_ULOGIC;
        RD5    : OUT STD_ULOGIC;
        RD4    : OUT STD_ULOGIC;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  
end component; 

component RAM8RA
  GENERIC (
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD7      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD6      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD5      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD4      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RDAD4_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_WRAD4_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC;
        RD6    : OUT STD_ULOGIC;
        RD5    : OUT STD_ULOGIC;
        RD4    : OUT STD_ULOGIC;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  
end component; 

component RAM8RF
  GENERIC (
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD7      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD6      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD5      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD4      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD4_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC;
        RD6    : OUT STD_ULOGIC;
        RD5    : OUT STD_ULOGIC;
        RD4    : OUT STD_ULOGIC;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  
end component; 

component RAM8RR
  GENERIC (
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD7      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD6      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD5      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD4      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD4_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC;
        RD6    : OUT STD_ULOGIC;
        RD5    : OUT STD_ULOGIC;
        RD4    : OUT STD_ULOGIC;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  
end component; 

component TBDLHS
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component TBHS
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component TF1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_T_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_T_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component TF1B
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_T_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_T_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
end component; 

component TRIBUFF
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
end component; 

component VCC
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True);

   port(
      Y                              :	out   STD_ULOGIC := '1');
end component; 

component XA1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component XA1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component XNOR2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component XO1
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component XO1A
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

component XOR2
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
end component; 

end COMPONENTS;

----------------------------------------------------------------
-- 
-- 
----------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;

library IEEE;
use IEEE.VITAL_Timing.all;
use IEEE.VITAL_Primitives.all;

package VTABLES is

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DF1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  S ),
    ( x,  x,  L,  x,  S ));

   CONSTANT DF1A_QN_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  H ),
    ( L,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  S ),
    ( x,  x,  L,  x,  S ));

   CONSTANT DFC1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  x,  L ),
    ( L,  H,  H,  L,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ));

   CONSTANT DFC1B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  H,  x,  L ));

   CONSTANT DFC1E_QN_tab : VitalStateTableType := (
    ( L,  H,  H,  H,  x,  L ),
    ( L,  x,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( x,  L,  x,  x,  x,  H ),
    ( x,  H,  x,  L,  x,  S ));

   CONSTANT DFE_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  L,  H,  H,  x,  L ),
    ( L,  x,  H,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   CONSTANT DFE3A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  H,  H,  x,  L ));

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ));

   CONSTANT DFM1B_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  L,  H,  x,  H ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  L,  x,  H,  x,  H ),
    ( L,  H,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  L,  H,  x,  H ),
    ( L,  x,  H,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   CONSTANT DFM3_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  x,  L ),
    ( L,  H,  H,  x,  H,  L,  x,  H ),
    ( L,  H,  x,  H,  H,  L,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  x,  L ),
    ( L,  x,  H,  L,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  x,  x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  x,  x,  H,  x,  L ));

   CONSTANT DFM4C_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  x,  L,  H,  x,  H ),
    ( H,  L,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  H,  H,  x,  H,  x,  L ),
    ( x,  L,  x,  H,  H,  H,  x,  L ));

   CONSTANT DFM6A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  H,  x,  L ));

   CONSTANT DFM7A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  x,  H,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  x,  H,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  L,  H,  x,  L ));

   CONSTANT DFME1A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( L,  L,  L,  x,  H,  x,  H,  x,  L ),
    ( L,  L,  x,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  H,  x,  x,  H,  x,  H ),
    ( L,  H,  H,  x,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  L,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  x,  L,  H,  x,  L ),
    ( L,  x,  L,  x,  H,  L,  H,  x,  L ),
    ( L,  x,  H,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  H,  x,  H,  L,  H,  x,  H ),
    ( L,  x,  x,  L,  L,  L,  H,  x,  L ),
    ( L,  x,  x,  H,  L,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  x,  x,  L,  x,  S ));

   CONSTANT DFP1_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  L,  x,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  H,  x,  x,  H ));

   CONSTANT DFP1B_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  S ),
    ( x,  x,  L,  x,  x,  H ),
    ( x,  x,  H,  L,  x,  S ));

   CONSTANT DFP1C_QN_tab : VitalStateTableType := (
    ( L,  L,  H,  L,  x,  H ),
    ( L,  H,  H,  x,  x,  L ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ));

   CONSTANT DFP1E_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  H,  H,  x,  L ));

   CONSTANT DFPC_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  H,  x,  H ),
    ( H,  H,  x,  L,  x,  x,  S ),
    ( H,  x,  x,  L,  L,  x,  S ),
    ( H,  x,  x,  H,  x,  x,  H ),
    ( x,  L,  L,  L,  H,  x,  L ));

   CONSTANT DL1_Q_tab : VitalStateTableType := (
    ( L,  H,  x,  L ),
    ( H,  H,  x,  H ),
    ( x,  L,  x,  S ));

   CONSTANT DL1A_QN_tab : VitalStateTableType := (
    ( L,  H,  x,  H ),
    ( H,  H,  x,  L ),
    ( x,  L,  x,  S ));

   CONSTANT DL1B_Q_tab : VitalStateTableType := (
    ( L,  L,  x,  L ),
    ( L,  H,  x,  H ),
    ( H,  x,  x,  S ));

   CONSTANT DL1C_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  H ),
    ( L,  H,  x,  L ),
    ( H,  x,  x,  S ));

   CONSTANT DL2A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  H,  x,  H,  x,  H ),
    ( H,  x,  L,  L,  x,  S ),
    ( H,  x,  H,  x,  x,  H ),
    ( x,  L,  L,  H,  x,  L ));

   CONSTANT DL2B_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  x,  x,  L ),
    ( L,  H,  H,  x,  x,  S ),
    ( L,  x,  L,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  H ),
    ( x,  H,  L,  L,  x,  H ));

   CONSTANT DL2C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  x,  H ),
    ( H,  H,  x,  L,  x,  S ),
    ( H,  x,  x,  H,  x,  H ),
    ( x,  L,  L,  L,  x,  L ));

   CONSTANT DL2D_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  x,  x,  L ),
    ( L,  H,  x,  L,  x,  S ),
    ( L,  x,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  H ),
    ( x,  H,  L,  H,  x,  H ));

   CONSTANT DLC_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  H,  H,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  L,  H,  x,  L ));

   CONSTANT DLC1_Q_tab : VitalStateTableType := (
    ( L,  H,  x,  x,  L ),
    ( H,  H,  L,  x,  H ),
    ( x,  L,  L,  x,  S ),
    ( x,  x,  H,  x,  L ));

   CONSTANT DLC1A_Q_tab : VitalStateTableType := (
    ( L,  L,  x,  x,  L ),
    ( L,  H,  L,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  x,  H,  x,  L ));

   CONSTANT DLC1F_QN_tab : VitalStateTableType := (
    ( L,  H,  H,  x,  L ),
    ( L,  x,  L,  x,  S ),
    ( H,  x,  x,  x,  H ),
    ( x,  L,  H,  x,  H ));

   CONSTANT DLC1G_QN_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( L,  x,  L,  x,  H ),
    ( H,  L,  x,  x,  S ),
    ( x,  H,  x,  x,  H ));

   CONSTANT DLCA_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  S ),
    ( x,  L,  L,  x,  L ));

   CONSTANT DLE_Q_tab : VitalStateTableType := (
    ( L,  H,  H,  x,  L ),
    ( H,  H,  H,  x,  H ),
    ( x,  L,  x,  x,  S ),
    ( x,  x,  L,  x,  S ));

   CONSTANT DLE1D_QN_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H ),
    ( L,  L,  H,  x,  L ),
    ( H,  x,  x,  x,  S ),
    ( x,  H,  x,  x,  S ));

   CONSTANT DLE2B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  H,  x,  x,  S ),
    ( x,  L,  L,  L,  x,  L ));

   CONSTANT DLE2C_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  x,  L ),
    ( L,  L,  H,  L,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  H,  x,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ));

   CONSTANT DLE3B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  L ),
    ( L,  L,  H,  x,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  H,  x,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  H ));

   CONSTANT DLE3C_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  H,  x,  L ),
    ( L,  L,  H,  x,  x,  H ),
    ( H,  x,  x,  H,  x,  S ),
    ( x,  H,  x,  H,  x,  S ),
    ( x,  x,  x,  L,  x,  H ));

   CONSTANT DLEC_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  L ),
    ( L,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  S ),
    ( x,  H,  x,  x,  S ));

   CONSTANT DLM_Q_tab : VitalStateTableType := (
    ( L,  L,  x,  H,  x,  L ),
    ( L,  x,  H,  H,  x,  L ),
    ( H,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  H,  x,  H ),
    ( x,  L,  L,  H,  x,  L ),
    ( x,  H,  L,  H,  x,  H ),
    ( x,  x,  x,  L,  x,  S ));

   CONSTANT DLM2_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  H,  H,  x,  H,  x,  H ),
    ( H,  H,  x,  H,  H,  x,  H ),
    ( H,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  H,  H,  x,  L ),
    ( x,  x,  L,  L,  H,  x,  L ));

   CONSTANT DLM2B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  S ),
    ( x,  L,  L,  L,  x,  x,  L ),
    ( x,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  x,  L ));

   CONSTANT DLM3_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  x,  x,  H,  H,  x,  L ),
    ( L,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( H,  H,  H,  H,  x,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( x,  L,  x,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  H,  x,  H,  x,  L,  H,  x,  H ),
    ( x,  H,  x,  x,  H,  L,  H,  x,  H ),
    ( x,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  x,  L,  x,  L,  H,  H,  x,  L ),
    ( x,  x,  H,  H,  L,  x,  H,  x,  H ),
    ( x,  x,  H,  x,  L,  H,  H,  x,  H ),
    ( x,  x,  x,  L,  L,  L,  H,  x,  L ),
    ( x,  x,  x,  H,  L,  L,  H,  x,  H ),
    ( x,  x,  x,  x,  x,  x,  L,  x,  S ));

   CONSTANT DLM3A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  L,  x,  x,  x,  L ),
    ( L,  L,  L,  x,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  L,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  H,  H,  x,  x,  x,  H ),
    ( L,  H,  H,  x,  x,  H,  x,  x,  H ),
    ( L,  H,  x,  H,  x,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  x,  L,  x,  L,  x,  L ),
    ( L,  x,  L,  x,  x,  H,  L,  x,  L ),
    ( L,  x,  H,  x,  H,  x,  L,  x,  H ),
    ( L,  x,  H,  x,  x,  H,  L,  x,  H ),
    ( L,  x,  x,  L,  L,  L,  x,  x,  L ),
    ( L,  x,  x,  L,  x,  L,  H,  x,  L ),
    ( L,  x,  x,  H,  H,  L,  x,  x,  H ),
    ( L,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  x,  x,  L,  L,  L,  x,  L ),
    ( L,  x,  x,  x,  H,  L,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  S ));

   CONSTANT DLM4_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  x,  x,  x,  H,  x,  H,  H,  x,  L ),
    ( L,  x,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( H,  H,  H,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  H,  x,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( x,  L,  x,  L,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  H,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( x,  H,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( x,  H,  x,  x,  x,  H,  L,  H,  x,  H ),
    ( x,  x,  L,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  x,  L,  x,  L,  L,  H,  H,  x,  L ),
    ( x,  x,  H,  H,  L,  L,  x,  H,  x,  H ),
    ( x,  x,  H,  x,  L,  L,  H,  H,  x,  H ),
    ( x,  x,  x,  L,  L,  L,  L,  H,  x,  L ),
    ( x,  x,  x,  H,  L,  L,  L,  H,  x,  H ),
    ( x,  x,  x,  x,  x,  x,  x,  L,  x,  S ));

   CONSTANT DLM4A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  L,  x,  x,  x,  x,  L ),
    ( L,  L,  L,  x,  x,  H,  x,  x,  x,  L ),
    ( L,  L,  L,  x,  x,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  L,  x,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  H,  H,  x,  x,  x,  x,  H ),
    ( L,  H,  H,  x,  x,  H,  x,  x,  x,  H ),
    ( L,  H,  H,  x,  x,  x,  H,  x,  x,  H ),
    ( L,  H,  x,  H,  x,  x,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  x,  L,  x,  x,  L,  x,  L ),
    ( L,  x,  L,  x,  x,  H,  x,  L,  x,  L ),
    ( L,  x,  L,  x,  x,  x,  H,  L,  x,  L ),
    ( L,  x,  H,  x,  H,  x,  x,  L,  x,  H ),
    ( L,  x,  H,  x,  x,  H,  x,  L,  x,  H ),
    ( L,  x,  H,  x,  x,  x,  H,  L,  x,  H ),
    ( L,  x,  x,  L,  L,  L,  L,  x,  x,  L ),
    ( L,  x,  x,  L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  x,  H,  H,  L,  L,  x,  x,  H ),
    ( L,  x,  x,  H,  x,  L,  L,  H,  x,  H ),
    ( L,  x,  x,  x,  L,  L,  L,  L,  x,  L ),
    ( L,  x,  x,  x,  H,  L,  L,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  S ));

   CONSTANT DLMA_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  x,  L ),
    ( L,  L,  x,  H,  x,  L ),
    ( L,  H,  H,  x,  x,  H ),
    ( L,  H,  x,  H,  x,  H ),
    ( L,  x,  L,  L,  x,  L ),
    ( L,  x,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  S ));

   CONSTANT DLME1A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  L ),
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  H,  H,  x,  x,  H ),
    ( L,  L,  H,  x,  H,  x,  H ),
    ( L,  L,  x,  L,  L,  x,  L ),
    ( L,  L,  x,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  H,  x,  x,  x,  x,  S ));

   CONSTANT DLP1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( H,  x,  H,  x,  H ),
    ( x,  L,  L,  x,  S ),
    ( x,  H,  x,  x,  H ));

   CONSTANT DLP1A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  L ),
    ( L,  H,  x,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  x,  H,  x,  H ));

   CONSTANT DLP1B_Q_tab : VitalStateTableType := (
    ( L,  H,  H,  x,  L ),
    ( H,  x,  H,  x,  H ),
    ( x,  L,  x,  x,  H ),
    ( x,  H,  L,  x,  S ));

   CONSTANT DLP1C_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( L,  H,  x,  x,  H ),
    ( H,  x,  H,  x,  S ),
    ( x,  x,  L,  x,  H ));

   CONSTANT DLP1D_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  H,  H,  x,  L ));

   CONSTANT DLP1E_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  L,  L,  x,  H ),
    ( H,  H,  x,  x,  S ),
    ( x,  L,  H,  x,  L ));

   CONSTANT TF1A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  H,  x,  H ),
    ( H,  L,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  H,  x,  L ),
    ( x,  L,  H,  H,  H,  x,  L ));


end VTABLES;

---- end of VITAL tables library ----
----- CELL AND2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND2 : entity is TRUE;
end AND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AND2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) AND (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND2_VITAL of AND2 is
   for VITAL_ACT
   end for;
end CFG_AND2_VITAL;


----- CELL AND2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND2A : entity is TRUE;
end AND2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AND2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) AND ((NOT A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND2A_VITAL of AND2A is
   for VITAL_ACT
   end for;
end CFG_AND2A_VITAL;


----- CELL AND2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND2B : entity is TRUE;
end AND2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AND2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) AND ((NOT A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND2B_VITAL of AND2B is
   for VITAL_ACT
   end for;
end CFG_AND2B_VITAL;


----- CELL AND3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND3 : entity is TRUE;
end AND3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AND3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) AND (A_ipd) AND (C_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND3_VITAL of AND3 is
   for VITAL_ACT
   end for;
end CFG_AND3_VITAL;


----- CELL AND3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND3A : entity is TRUE;
end AND3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AND3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) AND ((NOT A_ipd)) AND (C_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND3A_VITAL of AND3A is
   for VITAL_ACT
   end for;
end CFG_AND3A_VITAL;


----- CELL AND3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND3B : entity is TRUE;
end AND3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AND3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) AND ((NOT A_ipd)) AND (C_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND3B_VITAL of AND3B is
   for VITAL_ACT
   end for;
end CFG_AND3B_VITAL;


----- CELL AND3C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND3C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND3C : entity is TRUE;
end AND3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AND3C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND3C_VITAL of AND3C is
   for VITAL_ACT
   end for;
end CFG_AND3C_VITAL;


----- CELL AND4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND4 : entity is TRUE;
end AND4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AND4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) AND (A_ipd) AND (C_ipd) AND (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND4_VITAL of AND4 is
   for VITAL_ACT
   end for;
end CFG_AND4_VITAL;


----- CELL AND4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND4A : entity is TRUE;
end AND4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AND4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) AND ((NOT A_ipd)) AND (C_ipd) AND (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND4A_VITAL of AND4A is
   for VITAL_ACT
   end for;
end CFG_AND4A_VITAL;


----- CELL AND4B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND4B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND4B : entity is TRUE;
end AND4B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AND4B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) AND ((NOT A_ipd)) AND (C_ipd) AND (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 3 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND4B_VITAL of AND4B is
   for VITAL_ACT
   end for;
end CFG_AND4B_VITAL;


----- CELL AND4C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND4C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND4C : entity is TRUE;
end AND4C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AND4C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd)) AND (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND4C_VITAL of AND4C is
   for VITAL_ACT
   end for;
end CFG_AND4C_VITAL;


----- CELL AND4D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND4D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND4D : entity is TRUE;
end AND4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AND4D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd)) AND ((NOT D_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND4D_VITAL of AND4D is
   for VITAL_ACT
   end for;
end CFG_AND4D_VITAL;


----- CELL AND5B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AND5B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AND5B : entity is TRUE;
end AND5B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AND5B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((NOT B_ipd)) AND ((NOT A_ipd)) AND (C_ipd) AND (D_ipd) AND (E_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AND5B_VITAL of AND5B is
   for VITAL_ACT
   end for;
end CFG_AND5B_VITAL;


----- CELL AO1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO1 : entity is TRUE;
end AO1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR ((B_ipd) AND (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO1_VITAL of AO1 is
   for VITAL_ACT
   end for;
end CFG_AO1_VITAL;


----- CELL AO10 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO10 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO10 : entity is TRUE;
end AO10;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO10 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((E_ipd) OR (D_ipd)) AND ((C_ipd) OR ((B_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 4 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO10_VITAL of AO10 is
   for VITAL_ACT
   end for;
end CFG_AO10_VITAL;


----- CELL AO11 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO11 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO11 : entity is TRUE;
end AO11;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO11 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((C_ipd) AND ((B_ipd) OR (A_ipd))) OR ((B_ipd) AND (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO11_VITAL of AO11 is
   for VITAL_ACT
   end for;
end CFG_AO11_VITAL;


----- CELL AO1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO1A : entity is TRUE;
end AO1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR ((B_ipd) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO1A_VITAL of AO1A is
   for VITAL_ACT
   end for;
end CFG_AO1A_VITAL;


----- CELL AO1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO1B : entity is TRUE;
end AO1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) OR ((B_ipd) AND (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO1B_VITAL of AO1B is
   for VITAL_ACT
   end for;
end CFG_AO1B_VITAL;


----- CELL AO1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO1C : entity is TRUE;
end AO1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) OR ((B_ipd) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO1C_VITAL of AO1C is
   for VITAL_ACT
   end for;
end CFG_AO1C_VITAL;


----- CELL AO1D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO1D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO1D : entity is TRUE;
end AO1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO1D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR (((NOT B_ipd)) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO1D_VITAL of AO1D is
   for VITAL_ACT
   end for;
end CFG_AO1D_VITAL;


----- CELL AO1E -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO1E is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO1E : entity is TRUE;
end AO1E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO1E is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) OR (((NOT B_ipd)) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO1E_VITAL of AO1E is
   for VITAL_ACT
   end for;
end CFG_AO1E_VITAL;


----- CELL AO2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO2 : entity is TRUE;
end AO2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR ((B_ipd) AND (A_ipd)) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO2_VITAL of AO2 is
   for VITAL_ACT
   end for;
end CFG_AO2_VITAL;


----- CELL AO2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO2A : entity is TRUE;
end AO2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR ((B_ipd) AND ((NOT A_ipd))) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO2A_VITAL of AO2A is
   for VITAL_ACT
   end for;
end CFG_AO2A_VITAL;


----- CELL AO2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO2B : entity is TRUE;
end AO2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR (((NOT B_ipd)) AND ((NOT A_ipd))) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 3 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO2B_VITAL of AO2B is
   for VITAL_ACT
   end for;
end CFG_AO2B_VITAL;


----- CELL AO2C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO2C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO2C : entity is TRUE;
end AO2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO2C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) OR ((B_ipd) AND ((NOT A_ipd))) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO2C_VITAL of AO2C is
   for VITAL_ACT
   end for;
end CFG_AO2C_VITAL;


----- CELL AO2D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO2D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO2D : entity is TRUE;
end AO2D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO2D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((NOT C_ipd)) OR (((NOT B_ipd)) AND ((NOT A_ipd))) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO2D_VITAL of AO2D is
   for VITAL_ACT
   end for;
end CFG_AO2D_VITAL;


----- CELL AO2E -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO2E is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO2E : entity is TRUE;
end AO2E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO2E is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((NOT C_ipd)) OR (((NOT B_ipd)) AND ((NOT A_ipd))) OR ((NOT D_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO2E_VITAL of AO2E is
   for VITAL_ACT
   end for;
end CFG_AO2E_VITAL;


----- CELL AO3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO3 : entity is TRUE;
end AO3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (D_ipd) OR ((B_ipd) AND ((NOT A_ipd)) AND (C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO3_VITAL of AO3 is
   for VITAL_ACT
   end for;
end CFG_AO3_VITAL;


----- CELL AO3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO3A : entity is TRUE;
end AO3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (D_ipd) OR ((B_ipd) AND (A_ipd) AND (C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO3A_VITAL of AO3A is
   for VITAL_ACT
   end for;
end CFG_AO3A_VITAL;


----- CELL AO3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO3B : entity is TRUE;
end AO3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (D_ipd) OR (((NOT B_ipd)) AND ((NOT A_ipd)) AND (C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 3 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO3B_VITAL of AO3B is
   for VITAL_ACT
   end for;
end CFG_AO3B_VITAL;


----- CELL AO3C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO3C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO3C : entity is TRUE;
end AO3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO3C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (D_ipd) OR (((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO3C_VITAL of AO3C is
   for VITAL_ACT
   end for;
end CFG_AO3C_VITAL;


----- CELL AO4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO4A : entity is TRUE;
end AO4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of AO4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((C_ipd) AND (A_ipd) AND (D_ipd)) OR ((B_ipd) AND ((NOT A_ipd)) AND
         (C_ipd)) OR ((C_ipd) AND (B_ipd) AND (D_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO4A_VITAL of AO4A is
   for VITAL_ACT
   end for;
end CFG_AO4A_VITAL;


----- CELL AO5A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO5A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO5A : entity is TRUE;
end AO5A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of AO5A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((C_ipd) AND (A_ipd)) OR ((B_ipd) AND ((NOT A_ipd))) OR ((C_ipd) AND (B_ipd)) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO5A_VITAL of AO5A is
   for VITAL_ACT
   end for;
end CFG_AO5A_VITAL;


----- CELL AO6 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO6 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO6 : entity is TRUE;
end AO6;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO6 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((D_ipd) AND (C_ipd)) OR ((B_ipd) AND (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO6_VITAL of AO6 is
   for VITAL_ACT
   end for;
end CFG_AO6_VITAL;


----- CELL AO6A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO6A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO6A : entity is TRUE;
end AO6A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO6A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (((NOT D_ipd)) AND (C_ipd)) OR ((B_ipd) AND (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO6A_VITAL of AO6A is
   for VITAL_ACT
   end for;
end CFG_AO6A_VITAL;


----- CELL AO7 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO7 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO7 : entity is TRUE;
end AO7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO7 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (D_ipd) OR ((B_ipd) AND (A_ipd) AND (C_ipd)) OR (E_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 4 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO7_VITAL of AO7 is
   for VITAL_ACT
   end for;
end CFG_AO7_VITAL;


----- CELL AO8 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO8 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO8 : entity is TRUE;
end AO8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO8 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (((NOT D_ipd)) AND ((NOT C_ipd))) OR ((B_ipd) AND (A_ipd)) OR (E_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 4 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO8_VITAL of AO8 is
   for VITAL_ACT
   end for;
end CFG_AO8_VITAL;


----- CELL AO9 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AO9 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AO9 : entity is TRUE;
end AO9;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AO9 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR ((B_ipd) AND (A_ipd)) OR (D_ipd) OR (E_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 4 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AO9_VITAL of AO9 is
   for VITAL_ACT
   end for;
end CFG_AO9_VITAL;


----- CELL AOI1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI1 : entity is TRUE;
end AOI1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AOI1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((C_ipd) OR ((B_ipd) AND (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI1_VITAL of AOI1 is
   for VITAL_ACT
   end for;
end CFG_AOI1_VITAL;


----- CELL AOI1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI1A : entity is TRUE;
end AOI1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AOI1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((C_ipd) OR ((B_ipd) AND ((NOT A_ipd)))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI1A_VITAL of AOI1A is
   for VITAL_ACT
   end for;
end CFG_AOI1A_VITAL;


----- CELL AOI1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI1B : entity is TRUE;
end AOI1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AOI1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT C_ipd)) OR ((B_ipd) AND (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI1B_VITAL of AOI1B is
   for VITAL_ACT
   end for;
end CFG_AOI1B_VITAL;


----- CELL AOI1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI1C : entity is TRUE;
end AOI1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AOI1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((C_ipd) OR (((NOT B_ipd)) AND ((NOT A_ipd)))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI1C_VITAL of AOI1C is
   for VITAL_ACT
   end for;
end CFG_AOI1C_VITAL;


----- CELL AOI1D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI1D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI1D : entity is TRUE;
end AOI1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AOI1D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT C_ipd)) OR (((NOT B_ipd)) AND ((NOT A_ipd)))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI1D_VITAL of AOI1D is
   for VITAL_ACT
   end for;
end CFG_AOI1D_VITAL;


----- CELL AOI2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI2A : entity is TRUE;
end AOI2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AOI2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((C_ipd) OR ((B_ipd) AND ((NOT A_ipd))) OR (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI2A_VITAL of AOI2A is
   for VITAL_ACT
   end for;
end CFG_AOI2A_VITAL;


----- CELL AOI2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI2B : entity is TRUE;
end AOI2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AOI2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT C_ipd)) OR ((B_ipd) AND ((NOT A_ipd))) OR (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI2B_VITAL of AOI2B is
   for VITAL_ACT
   end for;
end CFG_AOI2B_VITAL;


----- CELL AOI3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI3A : entity is TRUE;
end AOI3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AOI3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((D_ipd) OR (A_ipd)) AND ((B_ipd) OR (A_ipd) OR (C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI3A_VITAL of AOI3A is
   for VITAL_ACT
   end for;
end CFG_AOI3A_VITAL;


----- CELL AOI4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI4 : entity is TRUE;
end AOI4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AOI4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((D_ipd) AND (C_ipd)) OR ((B_ipd) AND (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI4_VITAL of AOI4 is
   for VITAL_ACT
   end for;
end CFG_AOI4_VITAL;


----- CELL AOI4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AOI4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AOI4A : entity is TRUE;
end AOI4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AOI4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((D_ipd) AND ((NOT C_ipd))) OR ((B_ipd) AND (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AOI4A_VITAL of AOI4A is
   for VITAL_ACT
   end for;
end CFG_AOI4A_VITAL;


----- CELL AX1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AX1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AX1 : entity is TRUE;
end AX1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AX1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) XOR ((B_ipd) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AX1_VITAL of AX1 is
   for VITAL_ACT
   end for;
end CFG_AX1_VITAL;


----- CELL AX1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AX1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AX1A : entity is TRUE;
end AX1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AX1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((C_ipd) XOR ((B_ipd) AND ((NOT A_ipd)))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AX1A_VITAL of AX1A is
   for VITAL_ACT
   end for;
end CFG_AX1A_VITAL;


----- CELL AX1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AX1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AX1B : entity is TRUE;
end AX1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AX1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) XOR (((NOT B_ipd)) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AX1B_VITAL of AX1B is
   for VITAL_ACT
   end for;
end CFG_AX1B_VITAL;


----- CELL AX1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity AX1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of AX1C : entity is TRUE;
end AX1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of AX1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) XOR ((B_ipd) AND (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_AX1C_VITAL of AX1C is
   for VITAL_ACT
   end for;
end CFG_AX1C_VITAL;




----- CELL BBDLHS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BBDLHS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_GOUT_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_GIN_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_GOUT_noedge_negedge           :	VitalDelayType := 0.000 ns;
      tsetup_D_GOUT_noedge_negedge          :	VitalDelayType := 0.000 ns;
      thold_PAD_GIN_noedge_posedge          :	VitalDelayType := 0.000 ns;
      tsetup_PAD_GIN_noedge_posedge         :	VitalDelayType := 0.000 ns;
      tperiod_GIN_posedge            :	VitalDelayType := 0.000 ns;
      tperiod_GOUT_negedge           :	VitalDelayType := 0.000 ns;
      tpw_GIN_negedge                :	VitalDelayType := 0.000 ns;
      tpw_GOUT_posedge               :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_GIN                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_GOUT                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      GIN                            :	in    STD_ULOGIC;
      GOUT                           :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BBDLHS : entity is TRUE;
end BBDLHS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of BBDLHS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;


   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GIN_ipd	 : STD_ULOGIC := 'X';
   SIGNAL GOUT_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (GIN_ipd, GIN, tipd_GIN);
   VitalWireDelay (GOUT_ipd, GOUT, tipd_GOUT);
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, GIN_ipd, GOUT_ipd, PAD_ipd)


   -- timing check results
   VARIABLE Tviol_D_GOUT	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_GOUT	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PAD_GIN	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PAD_GIN	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_GOUT	: STD_ULOGIC := '0';
   VARIABLE PInfo_GOUT	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_GIN	: STD_ULOGIC := '0';
   VARIABLE PInfo_GIN	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_IQ : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 3) := (others => 'X');
   ALIAS IQ_zd : STD_LOGIC is Results(1);
   ALIAS Q_zd : STD_LOGIC is Results(2);
   ALIAS PAD_zd : STD_LOGIC is Results(3);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   -- State Table : DL1_Q_table Declaration
   CONSTANT DL1_Q_table : VitalStateTableType := (
    ( '0',  '1',  '-',  '0' ),
    ( '1',  '1',  '-',  '1' ),
    ( '-',  '0',  '-',  'S' ));

   -- State Table : DL1B_Q_table Declaration
   CONSTANT DL1B_Q_table : VitalStateTableType := (
    ( '0',  '0',  '-',  '0' ),
    ( '0',  '1',  '-',  '1' ),
    ( '1',  '-',  '-',  'S' ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_GOUT,
          TimingData              => Tmkr_D_GOUT,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => GOUT_ipd,
          RefSignalName          => "GOUT",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_GOUT_noedge_negedge,
          SetupLow                => tsetup_D_GOUT_noedge_negedge,
          HoldHigh                => thold_D_GOUT_noedge_negedge,
          HoldLow                 => thold_D_GOUT_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/BBDLHS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_PAD_GIN,
          TimingData              => Tmkr_PAD_GIN,
          TestSignal              => PAD_ipd,
          TestSignalName          => "PAD",
          TestDelay               => 0 ns,
          RefSignal               => GIN_ipd,
          RefSignalName          => "GIN",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_PAD_GIN_noedge_posedge,
          SetupLow                => tsetup_PAD_GIN_noedge_posedge,
          HoldHigh                => thold_PAD_GIN_noedge_posedge,
          HoldLow                 => thold_PAD_GIN_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/BBDLHS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GOUT,
          PeriodData              => PInfo_GOUT,
          TestSignal              => GOUT_ipd,
          TestSignalName          => "GOUT",
          TestDelay               => 0 ns,
          Period                  => tperiod_GOUT_negedge,
          PulseWidthHigh          => tpw_GOUT_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/BBDLHS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_GIN,
          PeriodData              => PInfo_GIN,
          TestSignal              => GIN_ipd,
          TestSignalName          => "GIN",
          TestDelay               => 0 ns,
          Period                  => tperiod_GIN_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_GIN_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/BBDLHS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_GOUT or Tviol_PAD_GIN or Pviol_GOUT or Pviol_GIN;
      VitalStateTable(
        Result => IQ_zd,
        PreviousDataIn => PrevData_IQ,
        StateTable => DL1_Q_table,
        DataIn => (
               D_ipd, GOUT_ipd));
      IQ_zd := Violation XOR IQ_zd;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DL1B_Q_table,
        DataIn => (
               GIN_ipd, PAD_ipd));
      Q_zd := Violation XOR Q_zd;
      PAD_zd := VitalBUFIF0 (data => IQ_zd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_PAD, TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE),
                 2 => (GOUT_ipd'last_event, VitalExtendToFillDelay(tpd_GOUT_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Q, TRUE),
                 1 => (GIN_ipd'last_event, tpd_GIN_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_BBDLHS_VITAL of BBDLHS is
   for VITAL_ACT
   end for;
end CFG_BBDLHS_VITAL;



----- CELL BBHS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BBHS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BBHS : entity is TRUE;
end BBHS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of BBHS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);
   ALIAS Y_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_PAD, TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_BBHS_VITAL of BBHS is
   for VITAL_ACT
   end for;
end CFG_BBHS_VITAL;


----- CELL BIBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BIBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BIBUF : entity is TRUE;
end BIBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of BIBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);
   ALIAS Y_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_PAD, TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_BIBUF_VITAL of BIBUF is
   for VITAL_ACT
   end for;
end CFG_BIBUF_VITAL;


----- CELL BUFA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFA : entity is TRUE;
end BUFA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of BUFA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_BUFA_VITAL of BUFA is
   for VITAL_ACT
   end for;
end CFG_BUFA_VITAL;


----- CELL BUFD -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFD is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFD : entity is TRUE;
end BUFD;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of BUFD is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_BUFD_VITAL of BUFD is
   for VITAL_ACT
   end for;
end CFG_BUFD_VITAL;


----- CELL BUFF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity BUFF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of BUFF : entity is TRUE;
end BUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of BUFF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_BUFF_VITAL of BUFF is
   for VITAL_ACT
   end for;
end CFG_BUFF_VITAL;


----- CELL CLKBIBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKBIBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	inout STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKBIBUF : entity is TRUE;
end CLKBIBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of CLKBIBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);
   ALIAS Y_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_PAD, TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CLKBIBUF_VITAL of CLKBIBUF is
   for VITAL_ACT
   end for;
end CFG_CLKBIBUF_VITAL;


----- CELL CLKBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKBUF : entity is TRUE;
end CLKBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of CLKBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CLKBUF_VITAL of CLKBUF is
   for VITAL_ACT
   end for;
end CFG_CLKBUF_VITAL;


----- CELL CLKINT -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CLKINT is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CLKINT : entity is TRUE;
end CLKINT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of CLKINT is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CLKINT_VITAL of CLKINT is
   for VITAL_ACT
   end for;
end CFG_CLKINT_VITAL;


----- CELL CM7 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CM7 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S11_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S10_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CM7 : entity is TRUE;
end CM7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CM7 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S10_ipd, S11_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   VARIABLE OR_Out, MUX1_Out, MUX2_Out : std_ulogic;

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      --Y_zd :=
      -- (((S11_ipd) OR (S10_ipd)) AND (((S0_ipd) AND (D3_ipd)) OR (((NOT
      --   S0_ipd)) AND (D2_ipd)))) OR (((NOT ((S11_ipd) OR (S10_ipd)))) AND
      --   (((S0_ipd) AND (D1_ipd)) OR (((NOT S0_ipd)) AND (D0_ipd))));
      OR_Out := VitalOR2(S10_ipd, S11_ipd);
      MUX1_Out := VitalMUX2(D1_ipd, D0_ipd, S0_ipd);
      MUX2_Out := VitalMUX2(D3_ipd, D2_ipd, S0_ipd);
      Y_zd := VitalMUX2(MUX2_Out, MUX1_Out, OR_Out);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S11_ipd'last_event, tpd_S11_Y, TRUE),
                 1 => (S10_ipd'last_event, tpd_S10_Y, TRUE),
                 2 => (S0_ipd'last_event, tpd_S0_Y, TRUE),
                 3 => (D3_ipd'last_event, tpd_D3_Y, TRUE),
                 4 => (D2_ipd'last_event, tpd_D2_Y, TRUE),
                 5 => (D1_ipd'last_event, tpd_D1_Y, TRUE),
                 6 => (D0_ipd'last_event, tpd_D0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CM7_VITAL of CM7 is
   for VITAL_ACT
   end for;
end CFG_CM7_VITAL;


----- CELL CM8 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CM8 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S11_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S10_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S01_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S00_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S00                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S01                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S10                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S11                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S00                            :	in    STD_ULOGIC;
      S01                            :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CM8 : entity is TRUE;
end CM8;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CM8 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S00_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S01_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S00_ipd, S00, tipd_S00);
   VitalWireDelay (S01_ipd, S01, tipd_S01);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S00_ipd, S01_ipd, S10_ipd, S11_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   VARIABLE AND_Out, OR_Out, MUX1_Out, MUX2_Out : std_ulogic;

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      --Y_zd :=
      -- (((S11_ipd) OR (S10_ipd)) AND (((S01_ipd) AND (S00_ipd) AND (D3_ipd))
      --   OR (((NOT ((S01_ipd) AND (S00_ipd)))) AND (D2_ipd)))) OR (((NOT
      --   ((S11_ipd) OR (S10_ipd)))) AND (((S01_ipd) AND (S00_ipd) AND
      --   (D1_ipd)) OR (((NOT ((S01_ipd) AND (S00_ipd)))) AND (D0_ipd))));
      AND_Out := VitalAND2(S00_ipd, S01_ipd);
      OR_Out := VitalOR2(S10_ipd, S11_ipd);
      MUX1_Out := VitalMUX2(D1_ipd, D0_ipd, AND_Out);
      MUX2_Out := VitalMUX2(D3_ipd, D2_ipd, AND_Out);
      Y_zd := VitalMUX2(MUX2_Out, MUX1_Out, OR_Out);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S11_ipd'last_event, tpd_S11_Y, TRUE),
                 1 => (S10_ipd'last_event, tpd_S10_Y, TRUE),
                 2 => (S01_ipd'last_event, tpd_S01_Y, TRUE),
                 3 => (S00_ipd'last_event, tpd_S00_Y, TRUE),
                 4 => (D3_ipd'last_event, tpd_D3_Y, TRUE),
                 5 => (D2_ipd'last_event, tpd_D2_Y, TRUE),
                 6 => (D1_ipd'last_event, tpd_D1_Y, TRUE),
                 7 => (D0_ipd'last_event, tpd_D0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CM8_VITAL of CM8 is
   for VITAL_ACT
   end for;
end CFG_CM8_VITAL;


----- CELL CS1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CS1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CS1 : entity is TRUE;
end CS1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CS1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   VARIABLE AND_Out, OR_Out : std_ulogic;

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      --Y_zd :=
      -- ((((B_ipd) AND (S_ipd)) OR (A_ipd)) AND (D_ipd)) OR ((C_ipd) AND
      --   ((NOT (((B_ipd) AND (S_ipd)) OR (A_ipd)))));
      AND_Out := VitalAND2(B_ipd, S_ipd);
      OR_Out := VitalOR2(A_ipd, AND_Out);
      Y_zd := VitalMUX2(D_ipd, C_ipd, OR_Out);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CS1_VITAL of CS1 is
   for VITAL_ACT
   end for;
end CFG_CS1_VITAL;


----- CELL CS2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CS2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CS2 : entity is TRUE;
end CS2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of CS2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   VARIABLE AND_Out, OR_Out : std_ulogic;

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      --Y_zd :=
      -- ((B_ipd) AND ((S_ipd) OR (A_ipd)) AND (D_ipd)) OR ((C_ipd) AND ((NOT
      --   ((B_ipd) AND ((S_ipd) OR (A_ipd))))));
      OR_Out := VitalOR2(A_ipd, S_ipd);
      AND_Out := VitalAND2(B_ipd, OR_Out);
      Y_zd := VitalMUX2(D_ipd, C_ipd, AND_Out);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CS2_VITAL of CS2 is
   for VITAL_ACT
   end for;
end CFG_CS2_VITAL;


----- CELL CY2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CY2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      A1                             :	in    STD_ULOGIC;
      B0                             :	in    STD_ULOGIC;
      B1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CY2A : entity is TRUE;
end CY2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of CY2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL A1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A0_ipd, A0, tipd_A0);
   VitalWireDelay (A1_ipd, A1, tipd_A1);
   VitalWireDelay (B0_ipd, B0, tipd_B0);
   VitalWireDelay (B1_ipd, B1, tipd_B1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A0_ipd, A1_ipd, B0_ipd, B1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((B0_ipd) AND (A0_ipd) AND (A1_ipd)) OR ((B1_ipd) AND (A1_ipd)) OR
         ((B0_ipd) AND (A0_ipd) AND (B1_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B1_ipd'last_event, tpd_B1_Y, TRUE),
                 1 => (B0_ipd'last_event, tpd_B0_Y, TRUE),
                 2 => (A1_ipd'last_event, tpd_A1_Y, TRUE),
                 3 => (A0_ipd'last_event, tpd_A0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CY2A_VITAL of CY2A is
   for VITAL_ACT
   end for;
end CFG_CY2A_VITAL;


----- CELL CY2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity CY2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      A1                             :	in    STD_ULOGIC;
      B0                             :	in    STD_ULOGIC;
      B1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of CY2B : entity is TRUE;
end CY2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of CY2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL A1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A0_ipd, A0, tipd_A0);
   VitalWireDelay (A1_ipd, A1, tipd_A1);
   VitalWireDelay (B0_ipd, B0, tipd_B0);
   VitalWireDelay (B1_ipd, B1, tipd_B1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A0_ipd, A1_ipd, B0_ipd, B1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((A1_ipd) AND ((B0_ipd) OR (A0_ipd))) OR ((B1_ipd) AND (A1_ipd)) OR
         ((B1_ipd) AND ((B0_ipd) OR (A0_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B1_ipd'last_event, tpd_B1_Y, TRUE),
                 1 => (B0_ipd'last_event, tpd_B0_Y, TRUE),
                 2 => (A1_ipd'last_event, tpd_A1_Y, TRUE),
                 3 => (A0_ipd'last_event, tpd_A0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_CY2B_VITAL of CY2B is
   for VITAL_ACT
   end for;
end CFG_CY2B_VITAL;


----- CELL DF1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1 : entity is TRUE;
end DF1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DF1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DF1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1_VITAL of DF1 is
   for VITAL_ACT
   end for;
end CFG_DF1_VITAL;


----- CELL DF1_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1_CC : entity is TRUE;
end DF1_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DF1_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DF1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1_CC_VITAL of DF1_CC is
   for VITAL_ACT
   end for;
end CFG_DF1_CC_VITAL;


----- CELL DF1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1A : entity is TRUE;
end DF1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DF1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DF1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DF1A_QN_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1A_VITAL of DF1A is
   for VITAL_ACT
   end for;
end CFG_DF1A_VITAL;


----- CELL DF1A_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1A_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1A_CC : entity is TRUE;
end DF1A_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DF1A_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DF1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DF1A_QN_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1A_CC_VITAL of DF1A_CC is
   for VITAL_ACT
   end for;
end CFG_DF1A_CC_VITAL;


----- CELL DF1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1B : entity is TRUE;
end DF1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DF1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1B_VITAL of DF1B is
   for VITAL_ACT
   end for;
end CFG_DF1B_VITAL;


----- CELL DF1B_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1B_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1B_CC : entity is TRUE;
end DF1B_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DF1B_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DF1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1B_CC_VITAL of DF1B_CC is
   for VITAL_ACT
   end for;
end CFG_DF1B_CC_VITAL;


----- CELL DF1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1C : entity is TRUE;
end DF1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DF1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DF1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DF1A_QN_tab,
        DataIn => (
               CLK_ipd, D_delayed, CLK_delayed));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1C_VITAL of DF1C is
   for VITAL_ACT
   end for;
end CFG_DF1C_VITAL;


----- CELL DF1C_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DF1C_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DF1C_CC : entity is TRUE;
end DF1C_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DF1C_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DF1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DF1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DF1A_QN_tab,
        DataIn => (
               CLK_ipd, D_delayed, CLK_delayed));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DF1C_CC_VITAL of DF1C_CC is
   for VITAL_ACT
   end for;
end CFG_DF1C_CC_VITAL;


----- CELL DFC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1 : entity is TRUE;
end DFC1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)


   CONSTANT DFC1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  x,  L ),
    ( L,  H,  H,  L,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1_VITAL of DFC1 is
   for VITAL_ACT
   end for;
end CFG_DFC1_VITAL;


----- CELL DFC1_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1_CC : entity is TRUE;
end DFC1_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  x,  L ),
    ( L,  H,  H,  L,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1_CC_VITAL of DFC1_CC is
   for VITAL_ACT
   end for;
end CFG_DFC1_CC_VITAL;


----- CELL DFC1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1A : entity is TRUE;
end DFC1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  x,  L ),
    ( L,  H,  H,  L,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, CLK_delayed, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1A_VITAL of DFC1A is
   for VITAL_ACT
   end for;
end CFG_DFC1A_VITAL;


----- CELL DFC1A_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1A_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1A_CC : entity is TRUE;
end DFC1A_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1A_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  x,  L ),
    ( L,  H,  H,  L,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, CLK_delayed, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1A_CC_VITAL of DFC1A_CC is
   for VITAL_ACT
   end for;
end CFG_DFC1A_CC_VITAL;


----- CELL DFC1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1B : entity is TRUE;
end DFC1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1B_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, D_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1B_VITAL of DFC1B is
   for VITAL_ACT
   end for;
end CFG_DFC1B_VITAL;


----- CELL DFC1B_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1B_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1B_CC : entity is TRUE;
end DFC1B_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1B_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1B_CC_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1B_CC_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, D_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1B_CC_VITAL of DFC1B_CC is
   for VITAL_ACT
   end for;
end CFG_DFC1B_CC_VITAL;


----- CELL DFC1D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1D : entity is TRUE;
end DFC1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1B_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, D_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1D_VITAL of DFC1D is
   for VITAL_ACT
   end for;
end CFG_DFC1D_VITAL;


----- CELL DFC1D_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1D_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1D_CC : entity is TRUE;
end DFC1D_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1D_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  L ));


   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFC1B_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, D_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1D_CC_VITAL of DFC1D_CC is
   for VITAL_ACT
   end for;
end CFG_DFC1D_CC_VITAL;


----- CELL DFC1E -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1E is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1E : entity is TRUE;
end DFC1E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1E is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1E_QN_tab : VitalStateTableType := (
    ( L,  H,  H,  H,  x,  L ),
    ( L,  x,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( x,  L,  x,  x,  x,  H ),
    ( x,  H,  x,  L,  x,  S ),
    ( x,  U,  x,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFC1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFC1E_QN_tab,
        DataIn => (
               CLK_delayed, CLR_ipd, D_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1E_VITAL of DFC1E is
   for VITAL_ACT
   end for;
end CFG_DFC1E_VITAL;


----- CELL DFC1G -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFC1G is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFC1G : entity is TRUE;
end DFC1G;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFC1G is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFC1E_QN_tab : VitalStateTableType := (
    ( L,  H,  H,  H,  x,  L ),
    ( L,  x,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( x,  L,  x,  x,  x,  H ),
    ( x,  H,  x,  L,  x,  S ),
    ( x,  U,  x,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFC1E_QN_tab,
        DataIn => (
               CLK_ipd, CLR_ipd, D_delayed, CLK_delayed));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFC1G_VITAL of DFC1G is
   for VITAL_ACT
   end for;
end CFG_DFC1G_VITAL;


----- CELL DFE -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE : entity is TRUE;
end DFE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  L,  H,  H,  x,  L ),
    ( L,  x,  H,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( E_ipd ) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE_Q_tab,
        DataIn => (
               CLK_delayed, Q_zd, D_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE_VITAL of DFE is
   for VITAL_ACT
   end for;
end CFG_DFE_VITAL;


----- CELL DFE_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE_CC : entity is TRUE;
end DFE_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  L,  H,  H,  x,  L ),
    ( L,  x,  H,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( E_ipd ) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE_Q_tab,
        DataIn => (
               CLK_delayed, Q_zd, D_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE_CC_VITAL of DFE_CC is
   for VITAL_ACT
   end for;
end CFG_DFE_CC_VITAL;


----- CELL DFE1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE1B : entity is TRUE;
end DFE1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT E_ipd)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_delayed, Q_zd, D_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE1B_VITAL of DFE1B is
   for VITAL_ACT
   end for;
end CFG_DFE1B_VITAL;


----- CELL DFE1B_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE1B_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE1B_CC : entity is TRUE;
end DFE1B_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE1B_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)


   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT E_ipd)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_delayed, Q_zd, D_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE1B_CC_VITAL of DFE1B_CC is
   for VITAL_ACT
   end for;
end CFG_DFE1B_CC_VITAL;


----- CELL DFE1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE1C : entity is TRUE;
end DFE1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT E_ipd)) /= '0' ,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_negedge,
          TimingData              => Tmkr_E_CLK_negedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_negedge,
          SetupLow                => tsetup_E_CLK_noedge_negedge,
          HoldHigh                => thold_E_CLK_noedge_negedge,
          HoldLow                 => thold_E_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_E_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_ipd, Q_zd, D_delayed, E_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE1C_VITAL of DFE1C is
   for VITAL_ACT
   end for;
end CFG_DFE1C_VITAL;


----- CELL DFE1C_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE1C_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE1C_CC : entity is TRUE;
end DFE1C_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE1C_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT E_ipd)) /= '0' ,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_negedge,
          TimingData              => Tmkr_E_CLK_negedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_negedge,
          SetupLow                => tsetup_E_CLK_noedge_negedge,
          HoldHigh                => thold_E_CLK_noedge_negedge,
          HoldLow                 => thold_E_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_E_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_ipd, Q_zd, D_delayed, E_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE1C_CC_VITAL of DFE1C_CC is
   for VITAL_ACT
   end for;
end CFG_DFE1C_CC_VITAL;


----- CELL DFE3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE3A : entity is TRUE;
end DFE3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  H,  H,  x,  L ),
    ( U,  x,  L,  x,  x,  x,  x,  L ));


   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(( CLR_ipd ) AND ( E_ipd )) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFE3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, Q_zd, D_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE3A_VITAL of DFE3A is
   for VITAL_ACT
   end for;
end CFG_DFE3A_VITAL;


----- CELL DFE3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE3B : entity is TRUE;
end DFE3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  H,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  H,  H,  x,  L ),
    ( U,  x,  L,  x,  x,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(( CLR_ipd ) AND ( E_ipd )) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_negedge,
          TimingData              => Tmkr_E_CLK_negedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_negedge,
          SetupLow                => tsetup_E_CLK_noedge_negedge,
          HoldHigh                => thold_E_CLK_noedge_negedge,
          HoldLow                 => thold_E_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_E_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, Q_zd, D_delayed, E_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE3B_VITAL of DFE3B is
   for VITAL_ACT
   end for;
end CFG_DFE3B_VITAL;


----- CELL DFE3C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE3C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE3C : entity is TRUE;
end DFE3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE3C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  L,  x,  x,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_E_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, Q_zd, D_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE3C_VITAL of DFE3C is
   for VITAL_ACT
   end for;
end CFG_DFE3C_VITAL;


----- CELL DFE3D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFE3D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFE3D : entity is TRUE;
end DFE3D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFE3D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  L,  x,  x,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE3D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_negedge,
          TimingData              => Tmkr_E_CLK_negedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_negedge,
          SetupLow                => tsetup_E_CLK_noedge_negedge,
          HoldHigh                => thold_E_CLK_noedge_negedge,
          HoldLow                 => thold_E_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE3D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFE3D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFE3D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFE3D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_E_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, Q_zd, D_delayed, E_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFE3D_VITAL of DFE3D is
   for VITAL_ACT
   end for;
end CFG_DFE3D_VITAL;


----- CELL DFEA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFEA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFEA : entity is TRUE;
end DFEA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFEA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  L,  H,  H,  x,  L ),
    ( L,  x,  H,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( E_ipd ) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFEA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_negedge,
          TimingData              => Tmkr_E_CLK_negedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_negedge,
          SetupLow                => tsetup_E_CLK_noedge_negedge,
          HoldHigh                => thold_E_CLK_noedge_negedge,
          HoldLow                 => thold_E_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFEA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFEA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_E_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE_Q_tab,
        DataIn => (
               CLK_ipd, Q_zd, D_delayed, E_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFEA_VITAL of DFEA is
   for VITAL_ACT
   end for;
end CFG_DFEA_VITAL;


----- CELL DFEA_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFEA_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFEA_CC : entity is TRUE;
end DFEA_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFEA_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  L,  H,  H,  x,  L ),
    ( L,  x,  H,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( E_ipd ) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFEA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_negedge,
          TimingData              => Tmkr_E_CLK_negedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_negedge,
          SetupLow                => tsetup_E_CLK_noedge_negedge,
          HoldHigh                => thold_E_CLK_noedge_negedge,
          HoldLow                 => thold_E_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFEA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFEA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Tviol_E_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE_Q_tab,
        DataIn => (
               CLK_ipd, Q_zd, D_delayed, E_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFEA_CC_VITAL of DFEA_CC is
   for VITAL_ACT
   end for;
end CFG_DFEA_CC_VITAL;


----- CELL DFM -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM : entity is TRUE;
end DFM;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_delayed, B_delayed, A_delayed, S_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM_VITAL of DFM is
   for VITAL_ACT
   end for;
end CFG_DFM_VITAL;


----- CELL DFM_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM_CC : entity is TRUE;
end DFM_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_delayed, B_delayed, A_delayed, S_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM_CC_VITAL of DFM_CC is
   for VITAL_ACT
   end for;
end CFG_DFM_CC_VITAL;


----- CELL DFM1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM1B : entity is TRUE;
end DFM1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM1B_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  L,  H,  x,  H ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  L,  x,  H,  x,  H ),
    ( L,  H,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  L,  H,  x,  H ),
    ( L,  x,  H,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFM1B_QN_tab,
        DataIn => (
               CLK_delayed, S_delayed, B_delayed, A_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM1B_VITAL of DFM1B is
   for VITAL_ACT
   end for;
end CFG_DFM1B_VITAL;


----- CELL DFM1B_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM1B_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM1B_CC : entity is TRUE;
end DFM1B_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM1B_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM1B_CC_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  L,  H,  x,  H ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  L,  x,  H,  x,  H ),
    ( L,  H,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  L,  H,  x,  H ),
    ( L,  x,  H,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFM1B_CC_QN_tab,
        DataIn => (
               CLK_delayed, S_delayed, B_delayed, A_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM1B_CC_VITAL of DFM1B_CC is
   for VITAL_ACT
   end for;
end CFG_DFM1B_CC_VITAL;


----- CELL DFM1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM1C : entity is TRUE;
end DFM1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM1B_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  L,  H,  x,  H ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  L,  x,  H,  x,  H ),
    ( L,  H,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  L,  H,  x,  H ),
    ( L,  x,  H,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_negedge,
          TimingData              => Tmkr_A_CLK_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_negedge,
          SetupLow                => tsetup_A_CLK_noedge_negedge,
          HoldHigh                => thold_A_CLK_noedge_negedge,
          HoldLow                 => thold_A_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_negedge,
          TimingData              => Tmkr_B_CLK_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_negedge,
          SetupLow                => tsetup_B_CLK_noedge_negedge,
          HoldHigh                => thold_B_CLK_noedge_negedge,
          HoldLow                 => thold_B_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_negedge,
          TimingData              => Tmkr_S_CLK_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_negedge,
          SetupLow                => tsetup_S_CLK_noedge_negedge,
          HoldHigh                => thold_S_CLK_noedge_negedge,
          HoldLow                 => thold_S_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_negedge or Tviol_B_CLK_negedge or Tviol_S_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFM1B_QN_tab,
        DataIn => (
               CLK_ipd, S_delayed, B_delayed, A_delayed, CLK_delayed));
      QN_zd := Violation XOR QN_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM1C_VITAL of DFM1C is
   for VITAL_ACT
   end for;
end CFG_DFM1C_VITAL;


----- CELL DFM1C_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM1C_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM1C_CC : entity is TRUE;
end DFM1C_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM1C_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM1B_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  L,  H,  x,  H ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  L,  x,  H,  x,  H ),
    ( L,  H,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  L,  H,  x,  H ),
    ( L,  x,  H,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_negedge,
          TimingData              => Tmkr_A_CLK_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_negedge,
          SetupLow                => tsetup_A_CLK_noedge_negedge,
          HoldHigh                => thold_A_CLK_noedge_negedge,
          HoldLow                 => thold_A_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_negedge,
          TimingData              => Tmkr_B_CLK_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_negedge,
          SetupLow                => tsetup_B_CLK_noedge_negedge,
          HoldHigh                => thold_B_CLK_noedge_negedge,
          HoldLow                 => thold_B_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_negedge,
          TimingData              => Tmkr_S_CLK_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_negedge,
          SetupLow                => tsetup_S_CLK_noedge_negedge,
          HoldHigh                => thold_S_CLK_noedge_negedge,
          HoldLow                 => thold_S_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM1C_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_negedge or Tviol_B_CLK_negedge or Tviol_S_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFM1B_QN_tab,
        DataIn => (
               CLK_ipd, S_delayed, B_delayed, A_delayed, CLK_delayed));
      QN_zd := Violation XOR QN_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM1C_CC_VITAL of DFM1C_CC is
   for VITAL_ACT
   end for;
end CFG_DFM1C_CC_VITAL;


----- CELL DFM3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM3 : entity is TRUE;
end DFM3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM3_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  x,  L ),
    ( L,  H,  H,  x,  H,  L,  x,  H ),
    ( L,  H,  x,  H,  H,  L,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  x,  L ),
    ( L,  x,  H,  L,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  x,  x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLR or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM3_Q_tab,
        DataIn => (
               CLK_delayed, B_delayed, A_delayed, S_delayed, CLK_ipd, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM3_VITAL of DFM3 is
   for VITAL_ACT
   end for;
end CFG_DFM3_VITAL;


----- CELL DFM3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM3B : entity is TRUE;
end DFM3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_negedge,
          TimingData              => Tmkr_A_CLK_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_negedge,
          SetupLow                => tsetup_A_CLK_noedge_negedge,
          HoldHigh                => thold_A_CLK_noedge_negedge,
          HoldLow                 => thold_A_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_negedge,
          TimingData              => Tmkr_B_CLK_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_negedge,
          SetupLow                => tsetup_B_CLK_noedge_negedge,
          HoldHigh                => thold_B_CLK_noedge_negedge,
          HoldLow                 => thold_B_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_negedge,
          TimingData              => Tmkr_S_CLK_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_negedge,
          SetupLow                => tsetup_S_CLK_noedge_negedge,
          HoldHigh                => thold_S_CLK_noedge_negedge,
          HoldLow                 => thold_S_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_negedge or Tviol_B_CLK_negedge or Tviol_S_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, B_delayed, A_delayed, S_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM3B_VITAL of DFM3B is
   for VITAL_ACT
   end for;
end CFG_DFM3B_VITAL;


----- CELL DFM3E -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM3E is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM3E : entity is TRUE;
end DFM3E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM3E is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM3_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  x,  L ),
    ( L,  H,  H,  x,  H,  L,  x,  H ),
    ( L,  H,  x,  H,  H,  L,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  x,  L ),
    ( L,  x,  H,  L,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  x,  x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_negedge,
          TimingData              => Tmkr_A_CLK_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_negedge,
          SetupLow                => tsetup_A_CLK_noedge_negedge,
          HoldHigh                => thold_A_CLK_noedge_negedge,
          HoldLow                 => thold_A_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_negedge,
          TimingData              => Tmkr_B_CLK_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_negedge,
          SetupLow                => tsetup_B_CLK_noedge_negedge,
          HoldHigh                => thold_B_CLK_noedge_negedge,
          HoldLow                 => thold_B_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_negedge,
          TimingData              => Tmkr_S_CLK_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_negedge,
          SetupLow                => tsetup_S_CLK_noedge_negedge,
          HoldHigh                => thold_S_CLK_noedge_negedge,
          HoldLow                 => thold_S_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM3E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFM3E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM3E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_negedge or Tviol_B_CLK_negedge or Tviol_S_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM3_Q_tab,
        DataIn => (
               CLK_ipd, B_delayed, A_delayed, S_delayed, CLK_delayed, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM3E_VITAL of DFM3E is
   for VITAL_ACT
   end for;
end CFG_DFM3E_VITAL;


----- CELL DFM4C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM4C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM4C : entity is TRUE;
end DFM4C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM4C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM4C_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  x,  L,  H,  x,  H ),
    ( H,  L,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  H,  H,  x,  H,  x,  L ),
    ( x,  L,  x,  H,  H,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM4C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM4C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM4C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM4C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM4C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM4C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFM4C_QN_tab,
        DataIn => (
               PRE_ipd, CLK_delayed, S_delayed, B_delayed, A_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM4C_VITAL of DFM4C is
   for VITAL_ACT
   end for;
end CFG_DFM4C_VITAL;


----- CELL DFM4D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM4D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM4D : entity is TRUE;
end DFM4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM4D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM4C_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  x,  L,  H,  x,  H ),
    ( H,  L,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  H,  H,  x,  H,  x,  L ),
    ( x,  L,  x,  H,  H,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_negedge,
          TimingData              => Tmkr_A_CLK_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_negedge,
          SetupLow                => tsetup_A_CLK_noedge_negedge,
          HoldHigh                => thold_A_CLK_noedge_negedge,
          HoldLow                 => thold_A_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM4D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_negedge,
          TimingData              => Tmkr_B_CLK_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_negedge,
          SetupLow                => tsetup_B_CLK_noedge_negedge,
          HoldHigh                => thold_B_CLK_noedge_negedge,
          HoldLow                 => thold_B_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM4D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_negedge,
          TimingData              => Tmkr_S_CLK_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_negedge,
          SetupLow                => tsetup_S_CLK_noedge_negedge,
          HoldHigh                => thold_S_CLK_noedge_negedge,
          HoldLow                 => thold_S_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM4D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM4D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM4D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM4D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_negedge or Pviol_PRE or Tviol_B_CLK_negedge or Tviol_S_CLK_negedge or Tviol_PRE_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFM4C_QN_tab,
        DataIn => (
               PRE_ipd, CLK_ipd, S_delayed, B_delayed, A_delayed, CLK_delayed));
      QN_zd := Violation XOR QN_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM4D_VITAL of DFM4D is
   for VITAL_ACT
   end for;
end CFG_DFM4D_VITAL;


----- CELL DFM6A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM6A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S1_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S1_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM6A : entity is TRUE;
end DFM6A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM6A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S1_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D0_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S1_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S1_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 8);
   VARIABLE D0_delayed : STD_ULOGIC := 'X';
   VARIABLE D1_delayed : STD_ULOGIC := 'X';
   VARIABLE D2_delayed : STD_ULOGIC := 'X';
   VARIABLE D3_delayed : STD_ULOGIC := 'X';
   VARIABLE S0_delayed : STD_ULOGIC := 'X';
   VARIABLE S1_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM6A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_CLK_posedge,
          TimingData              => Tmkr_D0_CLK_posedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_CLK_noedge_posedge,
          SetupLow                => tsetup_D0_CLK_noedge_posedge,
          HoldHigh                => thold_D0_CLK_noedge_posedge,
          HoldLow                 => thold_D0_CLK_noedge_posedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( S0_ipd ) OR ( S1_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_CLK_posedge,
          TimingData              => Tmkr_D1_CLK_posedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_CLK_noedge_posedge,
          SetupLow                => tsetup_D1_CLK_noedge_posedge,
          HoldHigh                => thold_D1_CLK_noedge_posedge,
          HoldLow                 => thold_D1_CLK_noedge_posedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( NOT S0_ipd ) OR ( S1_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_CLK_posedge,
          TimingData              => Tmkr_D2_CLK_posedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_CLK_noedge_posedge,
          SetupLow                => tsetup_D2_CLK_noedge_posedge,
          HoldHigh                => thold_D2_CLK_noedge_posedge,
          HoldLow                 => thold_D2_CLK_noedge_posedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( S0_ipd ) OR ( NOT S1_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_CLK_posedge,
          TimingData              => Tmkr_D3_CLK_posedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_CLK_noedge_posedge,
          SetupLow                => tsetup_D3_CLK_noedge_posedge,
          HoldHigh                => thold_D3_CLK_noedge_posedge,
          HoldLow                 => thold_D3_CLK_noedge_posedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( NOT S0_ipd ) OR ( NOT S1_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_CLK_posedge,
          TimingData              => Tmkr_S0_CLK_posedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_CLK_noedge_posedge,
          SetupLow                => tsetup_S0_CLK_noedge_posedge,
          HoldHigh                => thold_S0_CLK_noedge_posedge,
          HoldLow                 => thold_S0_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S1_CLK_posedge,
          TimingData              => Tmkr_S1_CLK_posedge,
          TestSignal              => S1_ipd,
          TestSignalName          => "S1",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S1_CLK_noedge_posedge,
          SetupLow                => tsetup_S1_CLK_noedge_posedge,
          HoldHigh                => thold_S1_CLK_noedge_posedge,
          HoldLow                 => thold_S1_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM6A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_CLK_posedge or Tviol_D3_CLK_posedge or Tviol_S1_CLK_posedge or Tviol_CLR_CLK_posedge or Tviol_D1_CLK_posedge or Tviol_D2_CLK_posedge or Tviol_S0_CLK_posedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM6A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, D3_delayed, D2_delayed, D1_delayed, D0_delayed, S1_delayed, S0_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D0_delayed := D0_ipd;
      D1_delayed := D1_ipd;
      D2_delayed := D2_ipd;
      D3_delayed := D3_ipd;
      S0_delayed := S0_ipd;
      S1_delayed := S1_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM6A_VITAL of DFM6A is
   for VITAL_ACT
   end for;
end CFG_DFM6A_VITAL;


----- CELL DFM6B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM6B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S1_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S1_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM6B : entity is TRUE;
end DFM6B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM6B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S1_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D0_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S1_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S1_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 8);
   VARIABLE D0_delayed : STD_ULOGIC := 'X';
   VARIABLE D1_delayed : STD_ULOGIC := 'X';
   VARIABLE D2_delayed : STD_ULOGIC := 'X';
   VARIABLE D3_delayed : STD_ULOGIC := 'X';
   VARIABLE S0_delayed : STD_ULOGIC := 'X';
   VARIABLE S1_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM6A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_CLK_negedge,
          TimingData              => Tmkr_D0_CLK_negedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_CLK_noedge_negedge,
          SetupLow                => tsetup_D0_CLK_noedge_negedge,
          HoldHigh                => thold_D0_CLK_noedge_negedge,
          HoldLow                 => thold_D0_CLK_noedge_negedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( S0_ipd ) OR ( S1_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_CLK_negedge,
          TimingData              => Tmkr_D1_CLK_negedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_CLK_noedge_negedge,
          SetupLow                => tsetup_D1_CLK_noedge_negedge,
          HoldHigh                => thold_D1_CLK_noedge_negedge,
          HoldLow                 => thold_D1_CLK_noedge_negedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( NOT S0_ipd ) OR ( S1_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_CLK_negedge,
          TimingData              => Tmkr_D2_CLK_negedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_CLK_noedge_negedge,
          SetupLow                => tsetup_D2_CLK_noedge_negedge,
          HoldHigh                => thold_D2_CLK_noedge_negedge,
          HoldLow                 => thold_D2_CLK_noedge_negedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( S0_ipd ) OR ( NOT S1_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_CLK_negedge,
          TimingData              => Tmkr_D3_CLK_negedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_CLK_noedge_negedge,
          SetupLow                => tsetup_D3_CLK_noedge_negedge,
          HoldHigh                => thold_D3_CLK_noedge_negedge,
          HoldLow                 => thold_D3_CLK_noedge_negedge,
          CheckEnabled            => 
                   TO_X01((NOT CLR_ipd) OR ( NOT S0_ipd ) OR ( NOT S1_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_CLK_negedge,
          TimingData              => Tmkr_S0_CLK_negedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_CLK_noedge_negedge,
          SetupLow                => tsetup_S0_CLK_noedge_negedge,
          HoldHigh                => thold_S0_CLK_noedge_negedge,
          HoldLow                 => thold_S0_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S1_CLK_negedge,
          TimingData              => Tmkr_S1_CLK_negedge,
          TestSignal              => S1_ipd,
          TestSignalName          => "S1",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S1_CLK_noedge_negedge,
          SetupLow                => tsetup_S1_CLK_noedge_negedge,
          HoldHigh                => thold_S1_CLK_noedge_negedge,
          HoldLow                 => thold_S1_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM6B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_CLK_negedge or Tviol_D1_CLK_negedge or Tviol_D2_CLK_negedge or Tviol_S0_CLK_negedge or Tviol_D3_CLK_negedge or Tviol_S1_CLK_negedge or Pviol_CLR or Tviol_CLR_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM6A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, D3_delayed, D2_delayed, D1_delayed, D0_delayed, S1_delayed, S0_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D0_delayed := D0_ipd;
      D1_delayed := D1_ipd;
      D2_delayed := D2_ipd;
      D3_delayed := D3_ipd;
      S0_delayed := S0_ipd;
      S1_delayed := S1_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM6B_VITAL of DFM6B is
   for VITAL_ACT
   end for;
end CFG_DFM6B_VITAL;


----- CELL DFM7A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM7A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      thold_S10_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S10_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_S11_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S11_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM7A : entity is TRUE;
end DFM7A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM7A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S10_ipd, S11_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D0_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S10_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S10_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S11_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S11_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 9);
   VARIABLE D0_delayed : STD_ULOGIC := 'X';
   VARIABLE D1_delayed : STD_ULOGIC := 'X';
   VARIABLE D2_delayed : STD_ULOGIC := 'X';
   VARIABLE D3_delayed : STD_ULOGIC := 'X';
   VARIABLE S0_delayed : STD_ULOGIC := 'X';
   VARIABLE S10_delayed : STD_ULOGIC := 'X';
   VARIABLE S11_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM7A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  x,  H,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  x,  H,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_CLK_posedge,
          TimingData              => Tmkr_D0_CLK_posedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_CLK_noedge_posedge,
          SetupLow                => tsetup_D0_CLK_noedge_posedge,
          HoldHigh                => thold_D0_CLK_noedge_posedge,
          HoldLow                 => thold_D0_CLK_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S0_ipd )
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_CLK_posedge,
          TimingData              => Tmkr_D1_CLK_posedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_CLK_noedge_posedge,
          SetupLow                => tsetup_D1_CLK_noedge_posedge,
          HoldHigh                => thold_D1_CLK_noedge_posedge,
          HoldLow                 => thold_D1_CLK_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT S0_ipd )
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_CLK_posedge,
          TimingData              => Tmkr_D2_CLK_posedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_CLK_noedge_posedge,
          SetupLow                => tsetup_D2_CLK_noedge_posedge,
          HoldHigh                => thold_D2_CLK_noedge_posedge,
          HoldLow                 => thold_D2_CLK_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S0_ipd )
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_CLK_posedge,
          TimingData              => Tmkr_D3_CLK_posedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_CLK_noedge_posedge,
          SetupLow                => tsetup_D3_CLK_noedge_posedge,
          HoldHigh                => thold_D3_CLK_noedge_posedge,
          HoldLow                 => thold_D3_CLK_noedge_posedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT S0_ipd )
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_CLK_posedge,
          TimingData              => Tmkr_S0_CLK_posedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_CLK_noedge_posedge,
          SetupLow                => tsetup_S0_CLK_noedge_posedge,
          HoldHigh                => thold_S0_CLK_noedge_posedge,
          HoldLow                 => thold_S0_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S10_CLK_posedge,
          TimingData              => Tmkr_S10_CLK_posedge,
          TestSignal              => S10_ipd,
          TestSignalName          => "S10",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S10_CLK_noedge_posedge,
          SetupLow                => tsetup_S10_CLK_noedge_posedge,
          HoldHigh                => thold_S10_CLK_noedge_posedge,
          HoldLow                 => thold_S10_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S11_CLK_posedge,
          TimingData              => Tmkr_S11_CLK_posedge,
          TestSignal              => S11_ipd,
          TestSignalName          => "S11",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S11_CLK_noedge_posedge,
          SetupLow                => tsetup_S11_CLK_noedge_posedge,
          HoldHigh                => thold_S11_CLK_noedge_posedge,
          HoldLow                 => thold_S11_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM7A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_CLK_posedge or Tviol_D3_CLK_posedge or Tviol_S11_CLK_posedge or Tviol_CLR_CLK_posedge or Tviol_D1_CLK_posedge or Tviol_D2_CLK_posedge or Tviol_S0_CLK_posedge or Pviol_CLR or Tviol_S10_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM7A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, D3_delayed, D2_delayed, D1_delayed, D0_delayed, S11_delayed, S10_delayed, S0_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D0_delayed := D0_ipd;
      D1_delayed := D1_ipd;
      D2_delayed := D2_ipd;
      D3_delayed := D3_ipd;
      S0_delayed := S0_ipd;
      S10_delayed := S10_ipd;
      S11_delayed := S11_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM7A_VITAL of DFM7A is
   for VITAL_ACT
   end for;
end CFG_DFM7A_VITAL;


----- CELL DFM7B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFM7B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D1_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D1_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D2_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D2_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_D3_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_D3_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S0_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tsetup_S0_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      thold_S10_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S10_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_S11_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      tsetup_S11_CLK_noedge_negedge                 :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFM7B : entity is TRUE;
end DFM7B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFM7B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S10_ipd, S11_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D0_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S10_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S10_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S11_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S11_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 9);
   VARIABLE D0_delayed : STD_ULOGIC := 'X';
   VARIABLE D1_delayed : STD_ULOGIC := 'X';
   VARIABLE D2_delayed : STD_ULOGIC := 'X';
   VARIABLE D3_delayed : STD_ULOGIC := 'X';
   VARIABLE S0_delayed : STD_ULOGIC := 'X';
   VARIABLE S10_delayed : STD_ULOGIC := 'X';
   VARIABLE S11_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM7A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  H,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  L,  H,  H,  x,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  H,  x,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( H,  L,  x,  H,  x,  x,  x,  H,  L,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  H,  L,  L,  x,  H,  x,  H ),
    ( H,  L,  x,  x,  H,  x,  L,  L,  H,  H,  x,  H ),
    ( H,  L,  x,  x,  x,  H,  L,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  L,  L,  x,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( x,  L,  L,  L,  x,  x,  x,  H,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  H,  x,  H,  H,  x,  L ),
    ( x,  L,  L,  x,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  L,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  L,  x,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  x,  L,  x,  L,  L,  H,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  L,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_CLK_negedge,
          TimingData              => Tmkr_D0_CLK_negedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_CLK_noedge_negedge,
          SetupLow                => tsetup_D0_CLK_noedge_negedge,
          HoldHigh                => thold_D0_CLK_noedge_negedge,
          HoldLow                 => thold_D0_CLK_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S0_ipd )
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_CLK_negedge,
          TimingData              => Tmkr_D1_CLK_negedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_CLK_noedge_negedge,
          SetupLow                => tsetup_D1_CLK_noedge_negedge,
          HoldHigh                => thold_D1_CLK_noedge_negedge,
          HoldLow                 => thold_D1_CLK_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT S0_ipd )
                              OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_CLK_negedge,
          TimingData              => Tmkr_D2_CLK_negedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_CLK_noedge_negedge,
          SetupLow                => tsetup_D2_CLK_noedge_negedge,
          HoldHigh                => thold_D2_CLK_noedge_negedge,
          HoldLow                 => thold_D2_CLK_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( S0_ipd )
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_CLK_negedge,
          TimingData              => Tmkr_D3_CLK_negedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_CLK_noedge_negedge,
          SetupLow                => tsetup_D3_CLK_noedge_negedge,
          HoldHigh                => thold_D3_CLK_noedge_negedge,
          HoldLow                 => thold_D3_CLK_noedge_negedge,
          CheckEnabled            => 
              TO_X01( (NOT CLR_ipd) OR ( NOT S0_ipd )
                              OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_CLK_negedge,
          TimingData              => Tmkr_S0_CLK_negedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_CLK_noedge_negedge,
          SetupLow                => tsetup_S0_CLK_noedge_negedge,
          HoldHigh                => thold_S0_CLK_noedge_negedge,
          HoldLow                 => thold_S0_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S10_CLK_negedge,
          TimingData              => Tmkr_S10_CLK_negedge,
          TestSignal              => S10_ipd,
          TestSignalName          => "S10",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S10_CLK_noedge_negedge,
          SetupLow                => tsetup_S10_CLK_noedge_negedge,
          HoldHigh                => thold_S10_CLK_noedge_negedge,
          HoldLow                 => thold_S10_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S11_CLK_negedge,
          TimingData              => Tmkr_S11_CLK_negedge,
          TestSignal              => S11_ipd,
          TestSignalName          => "S11",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S11_CLK_noedge_negedge,
          SetupLow                => tsetup_S11_CLK_noedge_negedge,
          HoldHigh                => thold_S11_CLK_noedge_negedge,
          HoldLow                 => thold_S11_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFM7B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_CLK_negedge or Tviol_D1_CLK_negedge or Tviol_D2_CLK_negedge or Tviol_S0_CLK_negedge or Tviol_S10_CLK_negedge or Tviol_D3_CLK_negedge or Pviol_CLR or Tviol_S11_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM7A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, D3_delayed, D2_delayed, D1_delayed, D0_delayed, S11_delayed, S10_delayed, S0_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D0_delayed := D0_ipd;
      D1_delayed := D1_ipd;
      D2_delayed := D2_ipd;
      D3_delayed := D3_ipd;
      S0_delayed := S0_ipd;
      S10_delayed := S10_ipd;
      S11_delayed := S11_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFM7B_VITAL of DFM7B is
   for VITAL_ACT
   end for;
end CFG_DFM7B_VITAL;


----- CELL DFMA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFMA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFMA : entity is TRUE;
end DFMA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFMA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_negedge,
          TimingData              => Tmkr_A_CLK_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_negedge,
          SetupLow                => tsetup_A_CLK_noedge_negedge,
          HoldHigh                => thold_A_CLK_noedge_negedge,
          HoldLow                 => thold_A_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_negedge,
          TimingData              => Tmkr_B_CLK_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_negedge,
          SetupLow                => tsetup_B_CLK_noedge_negedge,
          HoldHigh                => thold_B_CLK_noedge_negedge,
          HoldLow                 => thold_B_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_negedge,
          TimingData              => Tmkr_S_CLK_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_negedge,
          SetupLow                => tsetup_S_CLK_noedge_negedge,
          HoldHigh                => thold_S_CLK_noedge_negedge,
          HoldLow                 => thold_S_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_negedge or Tviol_B_CLK_negedge or Tviol_S_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_ipd, B_delayed, A_delayed, S_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFMA_VITAL of DFMA is
   for VITAL_ACT
   end for;
end CFG_DFMA_VITAL;


----- CELL DFMA_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFMA_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFMA_CC : entity is TRUE;
end DFMA_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFMA_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE1B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_negedge,
          TimingData              => Tmkr_A_CLK_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_negedge,
          SetupLow                => tsetup_A_CLK_noedge_negedge,
          HoldHigh                => thold_A_CLK_noedge_negedge,
          HoldLow                 => thold_A_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFMA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_negedge,
          TimingData              => Tmkr_B_CLK_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_negedge,
          SetupLow                => tsetup_B_CLK_noedge_negedge,
          HoldHigh                => thold_B_CLK_noedge_negedge,
          HoldLow                 => thold_B_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFMA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_negedge,
          TimingData              => Tmkr_S_CLK_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_negedge,
          SetupLow                => tsetup_S_CLK_noedge_negedge,
          HoldHigh                => thold_S_CLK_noedge_negedge,
          HoldLow                 => thold_S_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFMA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFMA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_negedge or Tviol_B_CLK_negedge or Tviol_S_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_ipd, B_delayed, A_delayed, S_delayed, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFMA_CC_VITAL of DFMA_CC is
   for VITAL_ACT
   end for;
end CFG_DFMA_CC_VITAL;


----- CELL DFMB -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFMB is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFMB : entity is TRUE;
end DFMB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFMB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFMB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFMB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFMB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFMB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFMB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFMB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLR or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, B_delayed, A_delayed, S_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFMB_VITAL of DFMB is
   for VITAL_ACT
   end for;
end CFG_DFMB_VITAL;


----- CELL DFME1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFME1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_A_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_B_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_B_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_E_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_E_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFME1A : entity is TRUE;
end DFME1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFME1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_A_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_E_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_E_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE A_delayed : STD_ULOGIC := 'X';
   VARIABLE B_delayed : STD_ULOGIC := 'X';
   VARIABLE S_delayed : STD_ULOGIC := 'X';
   VARIABLE E_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFME1A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( L,  L,  L,  x,  H,  x,  H,  x,  L ),
    ( L,  L,  x,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  H,  x,  x,  H,  x,  H ),
    ( L,  H,  H,  x,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  H,  L,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  L,  x,  L,  H,  x,  L ),
    ( L,  x,  L,  x,  H,  L,  H,  x,  L ),
    ( L,  x,  H,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  H,  x,  H,  L,  H,  x,  H ),
    ( L,  x,  x,  L,  L,  L,  H,  x,  L ),
    ( L,  x,  x,  H,  L,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  S ),
    ( x,  x,  x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_CLK_posedge,
          TimingData              => Tmkr_A_CLK_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_CLK_noedge_posedge,
          SetupLow                => tsetup_A_CLK_noedge_posedge,
          HoldHigh                => thold_A_CLK_noedge_posedge,
          HoldLow                 => thold_A_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(E_ipd OR S_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_CLK_posedge,
          TimingData              => Tmkr_B_CLK_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_CLK_noedge_posedge,
          SetupLow                => tsetup_B_CLK_noedge_posedge,
          HoldHigh                => thold_B_CLK_noedge_posedge,
          HoldLow                 => thold_B_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(E_ipd OR (NOT S_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_CLK_posedge,
          TimingData              => Tmkr_S_CLK_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_CLK_noedge_posedge,
          SetupLow                => tsetup_S_CLK_noedge_posedge,
          HoldHigh                => thold_S_CLK_noedge_posedge,
          HoldLow                 => thold_S_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(E_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_E_CLK_posedge,
          TimingData              => Tmkr_E_CLK_posedge,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_E_CLK_noedge_posedge,
          SetupLow                => tsetup_E_CLK_noedge_posedge,
          HoldHigh                => thold_E_CLK_noedge_posedge,
          HoldLow                 => thold_E_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_CLK_posedge or Tviol_S_CLK_posedge or Tviol_E_CLK_posedge or Tviol_B_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFME1A_Q_tab,
        DataIn => (
               CLK_delayed, Q_zd, B_delayed, A_delayed, S_delayed, E_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      A_delayed := A_ipd;
      B_delayed := B_ipd;
      S_delayed := S_ipd;
      E_delayed := E_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFME1A_VITAL of DFME1A is
   for VITAL_ACT
   end for;
end CFG_DFME1A_VITAL;


----- CELL DFP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1 : entity is TRUE;
end DFP1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  L,  x,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  H,  x,  x,  H ),
    ( x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, PRE_ipd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1_VITAL of DFP1 is
   for VITAL_ACT
   end for;
end CFG_DFP1_VITAL;


----- CELL DFP1_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1_CC : entity is TRUE;
end DFP1_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1_CC_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  L,  x,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  H,  x,  x,  H ),
    ( x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1_CC_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, PRE_ipd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1_CC_VITAL of DFP1_CC is
   for VITAL_ACT
   end for;
end CFG_DFP1_CC_VITAL;


----- CELL DFP1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1A : entity is TRUE;
end DFP1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  L,  x,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  H,  x,  x,  H ),
    ( x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, PRE_ipd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1A_VITAL of DFP1A is
   for VITAL_ACT
   end for;
end CFG_DFP1A_VITAL;


----- CELL DFP1A_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1A_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1A_CC : entity is TRUE;
end DFP1A_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1A_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  L,  x,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  H,  x,  x,  H ),
    ( x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1A_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, PRE_ipd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1A_CC_VITAL of DFP1A_CC is
   for VITAL_ACT
   end for;
end CFG_DFP1A_CC_VITAL;


----- CELL DFP1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1B : entity is TRUE;
end DFP1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1B_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  S ),
    ( x,  x,  L,  x,  x,  H ),
    ( x,  x,  H,  L,  x,  S ),
    ( x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1B_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, PRE_ipd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1B_VITAL of DFP1B is
   for VITAL_ACT
   end for;
end CFG_DFP1B_VITAL;


----- CELL DFP1B_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1B_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1B_CC : entity is TRUE;
end DFP1B_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1B_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1B_CC_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  S ),
    ( x,  x,  L,  x,  x,  H ),
    ( x,  x,  H,  L,  x,  S ),
    ( x,  x,  U,  x,  H,  H ));


   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1B_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1B_CC_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, PRE_ipd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1B_CC_VITAL of DFP1B_CC is
   for VITAL_ACT
   end for;
end CFG_DFP1B_CC_VITAL;


----- CELL DFP1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1C : entity is TRUE;
end DFP1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1C_QN_tab : VitalStateTableType := (
    ( L,  L,  H,  L,  x,  H ),
    ( L,  H,  H,  x,  x,  L ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFP1C_QN_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd, PRE_ipd));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1C_VITAL of DFP1C is
   for VITAL_ACT
   end for;
end CFG_DFP1C_VITAL;


----- CELL DFP1D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1D : entity is TRUE;
end DFP1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1B_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  S ),
    ( x,  x,  L,  x,  x,  H ),
    ( x,  x,  H,  L,  x,  S ),
    ( x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1B_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, PRE_ipd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1D_VITAL of DFP1D is
   for VITAL_ACT
   end for;
end CFG_DFP1D_VITAL;


----- CELL DFP1D_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1D_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1D_CC : entity is TRUE;
end DFP1D_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1D_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1B_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  H,  x,  L ),
    ( L,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  S ),
    ( x,  x,  L,  x,  x,  H ),
    ( x,  x,  H,  L,  x,  S ),
    ( x,  x,  U,  x,  H,  H ));


   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1D_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFP1B_Q_tab,
        DataIn => (
               CLK_ipd, D_delayed, PRE_ipd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1D_CC_VITAL of DFP1D_CC is
   for VITAL_ACT
   end for;
end CFG_DFP1D_CC_VITAL;


----- CELL DFP1E -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1E is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1E : entity is TRUE;
end DFP1E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1E is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1E_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  H,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Pviol_PRE or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFP1E_QN_tab,
        DataIn => (
               PRE_ipd, CLK_delayed, D_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1E_VITAL of DFP1E is
   for VITAL_ACT
   end for;
end CFG_DFP1E_VITAL;


----- CELL DFP1F -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1F is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1F : entity is TRUE;
end DFP1F;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1F is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1C_QN_tab : VitalStateTableType := (
    ( L,  L,  H,  L,  x,  H ),
    ( L,  H,  H,  x,  x,  L ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFP1C_QN_tab,
        DataIn => (
               CLK_ipd, D_delayed, CLK_delayed, PRE_ipd));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1F_VITAL of DFP1F is
   for VITAL_ACT
   end for;
end CFG_DFP1F_VITAL;


----- CELL DFP1G -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFP1G is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFP1G : entity is TRUE;
end DFP1G;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFP1G is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFP1E_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  L,  H,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_posedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFP1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFP1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFP1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DFP1E_QN_tab,
        DataIn => (
               PRE_ipd, CLK_ipd, D_delayed, CLK_delayed));
      QN_zd := Violation XOR QN_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFP1G_VITAL of DFP1G is
   for VITAL_ACT
   end for;
end CFG_DFP1G_VITAL;


----- CELL DFPC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFPC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFPC : entity is TRUE;
end DFPC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFPC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFPC_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  H,  x,  H ),
    ( H,  H,  x,  L,  x,  x,  S ),
    ( H,  x,  x,  L,  L,  x,  S ),
    ( H,  x,  x,  H,  x,  x,  H ),
    ( x,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  L,  L ),
    ( H,  x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFPC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFPC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFPC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFPC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_PRE or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFPC_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, D_delayed, PRE_ipd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 2 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFPC_VITAL of DFPC is
   for VITAL_ACT
   end for;
end CFG_DFPC_VITAL;


----- CELL DFPC_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFPC_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFPC_CC : entity is TRUE;
end DFPC_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFPC_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFPC_CC_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  H,  x,  H ),
    ( H,  H,  x,  L,  x,  x,  S ),
    ( H,  x,  x,  L,  L,  x,  S ),
    ( H,  x,  x,  H,  x,  x,  H ),
    ( x,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  L,  L ),
    ( H,  x,  x,  U,  x,  H,  H ));


   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFPC_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_posedge,
          TimingData              => Tmkr_PRE_CLK_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_posedge,
          Removal                 => thold_PRE_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFPC_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DFPC_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPC_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPC_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFPC_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Tviol_PRE_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_PRE or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFPC_CC_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, D_delayed, PRE_ipd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 2 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFPC_CC_VITAL of DFPC_CC is
   for VITAL_ACT
   end for;
end CFG_DFPC_CC_VITAL;


----- CELL DFPCA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFPCA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFPCA : entity is TRUE;
end DFPCA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFPCA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFPCA_tab : VitalStateTableType := (
    ( L,  x,  x,  H,  x,  x,  U ),
    ( L,  x,  x,  L,  x,  x,  L ),
    ( H,  L,  H,  x,  H,  x,  H ),
    ( H,  H,  x,  L,  x,  x,  S ),
    ( H,  x,  x,  L,  L,  x,  S ),
    ( H,  x,  x,  H,  x,  x,  H ),
    ( x,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  L,  x,  L,  L ),
    ( H,  x,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFPCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFPCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFPCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFPCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFPCA_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, D_delayed, PRE_ipd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 2 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFPCA_VITAL of DFPCA is
   for VITAL_ACT
   end for;
end CFG_DFPCA_VITAL;


----- CELL DFPCA_CC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DFPCA_CC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_PRE_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_PRE_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DFPCA_CC : entity is TRUE;
end DFPCA_CC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DFPCA_CC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFPCA_CC_tab : VitalStateTableType := (
    ( L,  x,  x,  H,  x,  x,  U ),
    ( L,  x,  x,  L,  x,  x,  L ),
    ( H,  L,  H,  x,  H,  x,  H ),
    ( H,  H,  x,  L,  x,  x,  S ),
    ( H,  x,  x,  L,  L,  x,  S ),
    ( H,  x,  x,  H,  x,  x,  H ),
    ( x,  L,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  L,  x,  L,  L ),
    ( H,  x,  x,  U,  x,  H,  H ));


   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_negedge,
          TimingData              => Tmkr_D_CLK_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_negedge,
          SetupLow                => tsetup_D_CLK_noedge_negedge,
          HoldHigh                => thold_D_CLK_noedge_negedge,
          HoldLow                 => thold_D_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFPCA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_CLK_negedge,
          TimingData              => Tmkr_PRE_CLK_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_CLK_negedge_negedge,
          Removal                 => thold_PRE_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFPCA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DFPCA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPCA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DFPCA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DFPCA_CC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_negedge or Pviol_PRE or Tviol_PRE_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFPCA_CC_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, D_delayed, PRE_ipd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 1 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 2 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DFPCA_CC_VITAL of DFPCA_CC is
   for VITAL_ACT
   end for;
end CFG_DFPCA_CC_VITAL;


----- CELL DL1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL1 : entity is TRUE;
end DL1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DL1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DL1_Q_tab,
        DataIn => (
               D_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL1_VITAL of DL1 is
   for VITAL_ACT
   end for;
end CFG_DL1_VITAL;


----- CELL DL1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL1A : entity is TRUE;
end DL1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DL1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Pviol_G;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DL1A_QN_tab,
        DataIn => (
               D_ipd, G_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL1A_VITAL of DL1A is
   for VITAL_ACT
   end for;
end CFG_DL1A_VITAL;


----- CELL DL1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL1B : entity is TRUE;
end DL1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DL1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DL1B_Q_tab,
        DataIn => (
               G_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL1B_VITAL of DL1B is
   for VITAL_ACT
   end for;
end CFG_DL1B_VITAL;


----- CELL DL1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL1C : entity is TRUE;
end DL1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DL1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Pviol_G;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DL1C_QN_tab,
        DataIn => (
               G_ipd, D_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL1C_VITAL of DL1C is
   for VITAL_ACT
   end for;
end CFG_DL1C_VITAL;


----- CELL DL2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL2A : entity is TRUE;
end DL2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DL2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DL2A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  H,  x,  H,  x,  H ),
    ( H,  x,  L,  L,  x,  S ),
    ( H,  x,  H,  x,  x,  H ),
    ( x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  L ),
    ( H,  x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_negedge,
          TimingData              => Tmkr_PRE_G_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_negedge_negedge,
          Removal                 => thold_PRE_G_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_negedge,
          TimingData              => Tmkr_CLR_G_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_negedge,
          Removal                 => thold_CLR_G_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or Tviol_CLR_G_negedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DL2A_Q_tab,
        DataIn => (
               CLR_ipd, D_ipd, PRE_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 3 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL2A_VITAL of DL2A is
   for VITAL_ACT
   end for;
end CFG_DL2A_VITAL;


----- CELL DL2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL2B : entity is TRUE;
end DL2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DL2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DL2B_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  x,  x,  L ),
    ( L,  H,  H,  x,  x,  S ),
    ( L,  x,  L,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  H ),
    ( x,  H,  L,  L,  x,  H ),
    ( U,  x,  x,  x,  H,  H ),
    ( L,  U,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(( (NOT PRE_ipd) ) OR ( CLR_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_posedge,
          TimingData              => Tmkr_PRE_G_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_posedge_posedge,
          Removal                 => thold_PRE_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01( ( CLR_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_negedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT PRE_ipd) ) OR ( CLR_ipd ) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TO_X01( ( CLR_ipd ) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Tviol_CLR_G_posedge or Pviol_PRE or Pviol_G or Pviol_CLR;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DL2B_QN_tab,
        DataIn => (
               CLR_ipd, PRE_ipd, G_ipd, D_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 3 => (CLR_ipd'last_event, tpd_CLR_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL2B_VITAL of DL2B is
   for VITAL_ACT
   end for;
end CFG_DL2B_VITAL;


----- CELL DL2C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL2C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL2C : entity is TRUE;
end DL2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DL2C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DL2C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  x,  H ),
    ( H,  H,  x,  L,  x,  S ),
    ( H,  x,  x,  H,  x,  H ),
    ( x,  L,  L,  L,  x,  L ),
    ( U,  x,  x,  x,  L,  L ),
    ( H,  x,  x,  U,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_posedge,
          TimingData              => Tmkr_PRE_G_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_negedge_posedge,
          Removal                 => thold_PRE_G_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DL2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(( PRE_ipd ) OR ( (NOT CLR_ipd) ) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01( (NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Tviol_CLR_G_posedge or Pviol_PRE or Pviol_G or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DL2C_Q_tab,
        DataIn => (
               CLR_ipd, G_ipd, D_ipd, PRE_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE),
                 3 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL2C_VITAL of DL2C is
   for VITAL_ACT
   end for;
end CFG_DL2C_VITAL;


----- CELL DL2D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DL2D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DL2D : entity is TRUE;
end DL2D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DL2D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DL2D_QN_tab : VitalStateTableType := (
    ( L,  L,  x,  x,  x,  L ),
    ( L,  H,  x,  L,  x,  S ),
    ( L,  x,  H,  H,  x,  L ),
    ( H,  x,  x,  x,  x,  H ),
    ( x,  H,  L,  H,  x,  H ),
    ( U,  x,  x,  x,  H,  H ),
    ( L,  U,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(( (NOT PRE_ipd) ) OR ( CLR_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_negedge,
          TimingData              => Tmkr_PRE_G_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_posedge_negedge,
          Removal                 => thold_PRE_G_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TO_X01( ( CLR_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_negedge,
          TimingData              => Tmkr_CLR_G_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_negedge_negedge,
          Removal                 => thold_CLR_G_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DL2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(( (NOT PRE_ipd) ) OR ( CLR_ipd ) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TO_X01( ( CLR_ipd ) ) /= '1',
          HeaderMsg               => InstancePath &"/DL2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DL2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or Tviol_CLR_G_negedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DL2D_QN_tab,
        DataIn => (
               CLR_ipd, PRE_ipd, D_ipd, G_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE),
                 3 => (CLR_ipd'last_event, tpd_CLR_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DL2D_VITAL of DL2D is
   for VITAL_ACT
   end for;
end CFG_DL2D_VITAL;


----- CELL DLC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLC : entity is TRUE;
end DLC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLC_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  H,  H,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  L,  H,  x,  L ),
    ( U,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_negedge,
          TimingData              => Tmkr_CLR_G_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_negedge,
          Removal                 => thold_CLR_G_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_CLR_G_negedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLC_Q_tab,
        DataIn => (
               CLR_ipd, D_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLC_VITAL of DLC is
   for VITAL_ACT
   end for;
end CFG_DLC_VITAL;


----- CELL DLC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLC1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLC1 : entity is TRUE;
end DLC1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLC1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLC1_Q_tab : VitalStateTableType := (
    ( L,  H,  x,  x,  L ),
    ( H,  H,  L,  x,  H ),
    ( x,  L,  L,  x,  S ),
    ( x,  x,  H,  x,  L ),
    ( x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_negedge,
          TimingData              => Tmkr_CLR_G_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_negedge_negedge,
          Removal                 => thold_CLR_G_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLC1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_CLR_G_negedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLC1_Q_tab,
        DataIn => (
               D_ipd, G_ipd, CLR_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLC1_VITAL of DLC1 is
   for VITAL_ACT
   end for;
end CFG_DLC1_VITAL;


----- CELL DLC1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLC1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLC1A : entity is TRUE;
end DLC1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLC1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLC1A_Q_tab : VitalStateTableType := (
    ( L,  L,  x,  x,  L ),
    ( L,  H,  L,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  x,  H,  x,  L ),
    ( x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_negedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLC1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_CLR_G_posedge or Pviol_G or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLC1A_Q_tab,
        DataIn => (
               G_ipd, D_ipd, CLR_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLC1A_VITAL of DLC1A is
   for VITAL_ACT
   end for;
end CFG_DLC1A_VITAL;


----- CELL DLC1F -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLC1F is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLC1F : entity is TRUE;
end DLC1F;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLC1F is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLC1F_QN_tab : VitalStateTableType := (
    ( L,  H,  H,  x,  L ),
    ( L,  x,  L,  x,  S ),
    ( H,  x,  x,  x,  H ),
    ( x,  L,  H,  x,  H ),
    ( U,  x,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLC1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_negedge,
          TimingData              => Tmkr_CLR_G_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_negedge_negedge,
          Removal                 => thold_CLR_G_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLC1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLC1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLC1F",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_CLR_G_negedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DLC1F_QN_tab,
        DataIn => (
               CLR_ipd, D_ipd, G_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE),
                 2 => (CLR_ipd'last_event, tpd_CLR_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLC1F_VITAL of DLC1F is
   for VITAL_ACT
   end for;
end CFG_DLC1F_VITAL;


----- CELL DLC1G -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLC1G is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLC1G : entity is TRUE;
end DLC1G;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLC1G is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLC1G_QN_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( L,  x,  L,  x,  H ),
    ( H,  L,  x,  x,  S ),
    ( x,  H,  x,  x,  H ),
    ( x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_negedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLC1G",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_CLR_G_posedge or Pviol_G or Pviol_CLR;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DLC1G_QN_tab,
        DataIn => (
               G_ipd, CLR_ipd, D_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE),
                 2 => (CLR_ipd'last_event, tpd_CLR_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLC1G_VITAL of DLC1G is
   for VITAL_ACT
   end for;
end CFG_DLC1G_VITAL;


----- CELL DLCA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLCA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLCA : entity is TRUE;
end DLCA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLCA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLCA_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  S ),
    ( x,  L,  L,  x,  L ),
    ( U,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLCA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_CLR_G_posedge or Pviol_G or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLCA_Q_tab,
        DataIn => (
               CLR_ipd, G_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLCA_VITAL of DLCA is
   for VITAL_ACT
   end for;
end CFG_DLCA_VITAL;


----- CELL DLE -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLE is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_E_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLE : entity is TRUE;
end DLE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLE is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_E_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLE_Q_tab : VitalStateTableType := (
    ( L,  H,  H,  x,  L ),
    ( H,  H,  H,  x,  H ),
    ( x,  L,  x,  x,  S ),
    ( x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(E_ipd) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_negedge,
          TimingData              => Tmkr_D_E_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_negedge,
          SetupLow                => tsetup_D_E_noedge_negedge,
          HoldHigh                => thold_D_E_noedge_negedge,
          HoldLow                 => thold_D_E_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(G_ipd) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_E_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(G_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(E_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLE",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_D_E_negedge or Pviol_E or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLE_Q_tab,
        DataIn => (
               D_ipd, G_ipd, E_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLE_VITAL of DLE is
   for VITAL_ACT
   end for;
end CFG_DLE_VITAL;


----- CELL DLE1D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLE1D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLE1D : entity is TRUE;
end DLE1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLE1D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLE1D_QN_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H ),
    ( L,  L,  H,  x,  L ),
    ( H,  x,  x,  x,  S ),
    ( x,  H,  x,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(NOT E_ipd) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_posedge,
          TimingData              => Tmkr_D_E_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_posedge,
          SetupLow                => tsetup_D_E_noedge_posedge,
          HoldHigh                => thold_D_E_noedge_posedge,
          HoldLow                 => thold_D_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(NOT G_ipd) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TO_X01(NOT G_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLE1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(NOT E_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLE1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Pviol_E or Tviol_D_E_posedge or Pviol_G;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DLE1D_QN_tab,
        DataIn => (
               G_ipd, E_ipd, D_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (E_ipd'last_event, tpd_E_QN, TRUE),
                 2 => (G_ipd'last_event, tpd_G_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLE1D_VITAL of DLE1D is
   for VITAL_ACT
   end for;
end CFG_DLE1D_VITAL;


----- CELL DLE2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLE2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_CLR_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_CLR_E_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLE2B : entity is TRUE;
end DLE2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLE2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLE2B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  S ),
    ( H,  x,  H,  x,  x,  S ),
    ( x,  L,  L,  L,  x,  L ),
    ( U,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_posedge,
          TimingData              => Tmkr_D_E_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_posedge,
          SetupLow                => tsetup_D_E_noedge_posedge,
          HoldHigh                => thold_D_E_noedge_posedge,
          HoldLow                 => thold_D_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd) AND (NOT G_ipd)) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_E_posedge,
          TimingData              => Tmkr_CLR_E_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_E_posedge_posedge,
          Removal                 => thold_CLR_E_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            =>
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd) AND (NOT G_ipd)) /= '0',
          HeaderMsg               => InstancePath &"/DLE2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01((CLR_ipd) AND (NOT E_ipd)) /= '0',
          HeaderMsg               => InstancePath &"/DLE2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLE2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_CLR_G_posedge or Pviol_E or Tviol_D_E_posedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLE2B_Q_tab,
        DataIn => (
               CLR_ipd, G_ipd, E_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 3 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLE2B_VITAL of DLE2B is
   for VITAL_ACT
   end for;
end CFG_DLE2B_VITAL;


----- CELL DLE2C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLE2C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_CLR_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_CLR_E_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLE2C : entity is TRUE;
end DLE2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLE2C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLE2C_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  x,  L ),
    ( L,  L,  H,  L,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  H,  x,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  U,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd OR E_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_posedge,
          TimingData              => Tmkr_D_E_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_posedge,
          SetupLow                => tsetup_D_E_noedge_posedge,
          HoldHigh                => thold_D_E_noedge_posedge,
          HoldLow                 => thold_D_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd OR G_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_negedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_E_posedge,
          TimingData              => Tmkr_CLR_E_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_E_negedge_posedge,
          Removal                 => thold_CLR_E_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd OR G_ipd) /= '1',
          HeaderMsg               => InstancePath &"/DLE2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd OR E_ipd) /= '1',
          HeaderMsg               => InstancePath &"/DLE2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLE2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_CLR_G_posedge or Pviol_E or Tviol_D_E_posedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLE2C_Q_tab,
        DataIn => (
               G_ipd, E_ipd, D_ipd, CLR_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 3 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLE2C_VITAL of DLE2C is
   for VITAL_ACT
   end for;
end CFG_DLE2C_VITAL;


----- CELL DLE3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLE3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_PRE_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_PRE_E_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLE3B : entity is TRUE;
end DLE3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLE3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLE3B_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  L ),
    ( L,  L,  H,  x,  x,  H ),
    ( H,  x,  x,  L,  x,  S ),
    ( x,  H,  x,  L,  x,  S ),
    ( x,  x,  x,  H,  x,  H ),
    ( x,  x,  x,  U,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd OR E_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_posedge,
          TimingData              => Tmkr_D_E_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_posedge,
          SetupLow                => tsetup_D_E_noedge_posedge,
          HoldHigh                => thold_D_E_noedge_posedge,
          HoldLow                 => thold_D_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd OR G_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_posedge,
          TimingData              => Tmkr_PRE_G_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_negedge_posedge,
          Removal                 => thold_PRE_G_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_E_posedge,
          TimingData              => Tmkr_PRE_E_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_E_negedge_posedge,
          Removal                 => thold_PRE_E_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd OR G_ipd) /= '1',
          HeaderMsg               => InstancePath &"/DLE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd OR E_ipd) /= '1',
          HeaderMsg               => InstancePath &"/DLE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLE3B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_E or Pviol_PRE or Tviol_D_E_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLE3B_Q_tab,
        DataIn => (
               G_ipd, E_ipd, D_ipd, PRE_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 3 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLE3B_VITAL of DLE3B is
   for VITAL_ACT
   end for;
end CFG_DLE3B_VITAL;


----- CELL DLE3C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLE3C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_PRE_E_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      trecovery_PRE_E_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLE3C : entity is TRUE;
end DLE3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLE3C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLE3C_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  H,  x,  L ),
    ( L,  L,  H,  x,  x,  H ),
    ( H,  x,  x,  H,  x,  S ),
    ( x,  H,  x,  H,  x,  S ),
    ( x,  x,  x,  L,  x,  H ),
    ( x,  x,  x,  U,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) OR E_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_posedge,
          TimingData              => Tmkr_D_E_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_posedge,
          SetupLow                => tsetup_D_E_noedge_posedge,
          HoldHigh                => thold_D_E_noedge_posedge,
          HoldLow                 => thold_D_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) OR G_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_posedge,
          TimingData              => Tmkr_PRE_G_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_posedge_posedge,
          Removal                 => thold_PRE_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_E_posedge,
          TimingData              => Tmkr_PRE_E_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_E_posedge_posedge,
          Removal                 => thold_PRE_E_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) OR G_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) OR E_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLE3C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_E or Pviol_PRE or Tviol_D_E_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLE3C_Q_tab,
        DataIn => (
               G_ipd, E_ipd, D_ipd, PRE_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 3 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLE3C_VITAL of DLE3C is
   for VITAL_ACT
   end for;
end CFG_DLE3C_VITAL;


----- CELL DLEA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLEA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLEA : entity is TRUE;
end DLEA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLEA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DF1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  S ),
    ( x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_posedge,
          TimingData              => Tmkr_D_E_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_posedge,
          SetupLow                => tsetup_D_E_noedge_posedge,
          HoldHigh                => thold_D_E_noedge_posedge,
          HoldLow                 => thold_D_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(G_ipd) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLEA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(NOT E_ipd) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLEA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TO_X01(G_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLEA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(NOT E_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLEA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_E_posedge or Tviol_D_G_negedge or Pviol_E or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               E_ipd, D_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLEA_VITAL of DLEA is
   for VITAL_ACT
   end for;
end CFG_DLEA_VITAL;


----- CELL DLEB -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLEB is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_E_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLEB : entity is TRUE;
end DLEB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLEB is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_E_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DF1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( L,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  S ),
    ( x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_negedge,
          TimingData              => Tmkr_D_E_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_negedge,
          SetupLow                => tsetup_D_E_noedge_negedge,
          HoldHigh                => thold_D_E_noedge_negedge,
          HoldLow                 => thold_D_E_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(NOT G_ipd) /= '0',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLEB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(E_ipd) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLEB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_E_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(NOT G_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLEB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(E_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLEB",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_E_negedge or Pviol_E or Tviol_D_G_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               G_ipd, D_ipd, E_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLEB_VITAL of DLEB is
   for VITAL_ACT
   end for;
end CFG_DLEB_VITAL;


----- CELL DLEC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLEC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_D_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLEC : entity is TRUE;
end DLEC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLEC is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLEC_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  L ),
    ( L,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  S ),
    ( x,  H,  x,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(NOT E_ipd) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLEC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D_E_posedge,
          TimingData              => Tmkr_D_E_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_E_noedge_posedge,
          SetupLow                => tsetup_D_E_noedge_posedge,
          HoldHigh                => thold_D_E_noedge_posedge,
          HoldLow                 => thold_D_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(NOT G_ipd) /= '0',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLEC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TO_X01(NOT G_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLEC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(NOT E_ipd) /= '0',
          HeaderMsg               => InstancePath &"/DLEC",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Pviol_E or Tviol_D_E_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLEC_Q_tab,
        DataIn => (
               G_ipd, E_ipd, D_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 2 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLEC_VITAL of DLEC is
   for VITAL_ACT
   end for;
end CFG_DLEC_VITAL;


----- CELL DLM -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM : entity is TRUE;
end DLM;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_A_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM_Q_tab : VitalStateTableType := (
    ( L,  L,  x,  H,  x,  L ),
    ( L,  x,  H,  H,  x,  L ),
    ( H,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  H,  x,  H ),
    ( x,  L,  L,  H,  x,  L ),
    ( x,  H,  L,  H,  x,  H ),
    ( x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_G_negedge,
          TimingData              => Tmkr_A_G_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_G_noedge_negedge,
          SetupLow                => tsetup_A_G_noedge_negedge,
          HoldHigh                => thold_A_G_noedge_negedge,
          HoldLow                 => thold_A_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_G_negedge,
          TimingData              => Tmkr_B_G_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_G_noedge_negedge,
          SetupLow                => tsetup_B_G_noedge_negedge,
          HoldHigh                => thold_B_G_noedge_negedge,
          HoldLow                 => thold_B_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_G_negedge,
          TimingData              => Tmkr_S_G_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_G_noedge_negedge,
          SetupLow                => tsetup_S_G_noedge_negedge,
          HoldHigh                => thold_S_G_noedge_negedge,
          HoldLow                 => thold_S_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_G_negedge or Tviol_B_G_negedge or Tviol_S_G_negedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM_Q_tab,
        DataIn => (
               B_ipd, A_ipd, S_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE),
                 3 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM_VITAL of DLM is
   for VITAL_ACT
   end for;
end CFG_DLM_VITAL;


----- CELL DLM2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_A_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_B                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM2 : entity is TRUE;
end DLM2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_A_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM2_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  H,  H,  x,  H,  x,  H ),
    ( H,  H,  x,  H,  H,  x,  H ),
    ( H,  x,  H,  L,  H,  x,  H ),
    ( H,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  H,  H,  x,  L ),
    ( x,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_G_negedge,
          TimingData              => Tmkr_A_G_negedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_G_noedge_negedge,
          SetupLow                => tsetup_A_G_noedge_negedge,
          HoldHigh                => thold_A_G_noedge_negedge,
          HoldLow                 => thold_A_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM2",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_G_negedge,
          TimingData              => Tmkr_B_G_negedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_G_noedge_negedge,
          SetupLow                => tsetup_B_G_noedge_negedge,
          HoldHigh                => thold_B_G_noedge_negedge,
          HoldLow                 => thold_B_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM2",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_G_negedge,
          TimingData              => Tmkr_S_G_negedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_G_noedge_negedge,
          SetupLow                => tsetup_S_G_noedge_negedge,
          HoldHigh                => thold_S_G_noedge_negedge,
          HoldLow                 => thold_S_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM2",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_negedge,
          TimingData              => Tmkr_CLR_G_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_negedge,
          Removal                 => thold_CLR_G_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM2",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLM2",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM2",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_G_negedge or Tviol_B_G_negedge or Tviol_S_G_negedge or Pviol_CLR or Tviol_CLR_G_negedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM2_Q_tab,
        DataIn => (
               CLR_ipd, B_ipd, A_ipd, S_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE),
                 3 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 4 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM2_VITAL of DLM2 is
   for VITAL_ACT
   end for;
end CFG_DLM2_VITAL;


----- CELL DLM2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_CLR_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_A_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_CLR_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_CLR_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_B                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM2B : entity is TRUE;
end DLM2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, G_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_A_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM2B_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  x,  H ),
    ( H,  L,  H,  x,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  S ),
    ( x,  L,  L,  L,  x,  x,  L ),
    ( x,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  x,  L ),
    ( U,  x,  x,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_G_posedge,
          TimingData              => Tmkr_A_G_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_G_noedge_posedge,
          SetupLow                => tsetup_A_G_noedge_posedge,
          HoldHigh                => thold_A_G_noedge_posedge,
          HoldLow                 => thold_A_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_G_posedge,
          TimingData              => Tmkr_B_G_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_G_noedge_posedge,
          SetupLow                => tsetup_B_G_noedge_posedge,
          HoldHigh                => thold_B_G_noedge_posedge,
          HoldLow                 => thold_B_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd ) OR (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_G_posedge,
          TimingData              => Tmkr_S_G_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_G_noedge_posedge,
          SetupLow                => tsetup_S_G_noedge_posedge,
          HoldHigh                => thold_S_G_noedge_posedge,
          HoldLow                 => thold_S_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_G_posedge,
          TimingData              => Tmkr_CLR_G_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_G_posedge_posedge,
          Removal                 => thold_CLR_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLM2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_G_posedge or Tviol_B_G_posedge or Tviol_CLR_G_posedge or Tviol_S_G_posedge or Pviol_CLR or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM2B_Q_tab,
        DataIn => (
               CLR_ipd, G_ipd, B_ipd, A_ipd, S_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE),
                 3 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 4 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM2B_VITAL of DLM2B is
   for VITAL_ACT
   end for;
end CFG_DLM2B_VITAL;


----- CELL DLM3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S1_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S1_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM3 : entity is TRUE;
end DLM3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S1_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D0_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S1_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S1_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM3_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  x,  x,  H,  H,  x,  L ),
    ( L,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( H,  H,  H,  H,  x,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( x,  L,  x,  L,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  H,  x,  H,  x,  L,  H,  x,  H ),
    ( x,  H,  x,  x,  H,  L,  H,  x,  H ),
    ( x,  x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  x,  L,  x,  L,  H,  H,  x,  L ),
    ( x,  x,  H,  H,  L,  x,  H,  x,  H ),
    ( x,  x,  H,  x,  L,  H,  H,  x,  H ),
    ( x,  x,  x,  L,  L,  L,  H,  x,  L ),
    ( x,  x,  x,  H,  L,  L,  H,  x,  H ),
    ( x,  x,  x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_G_negedge,
          TimingData              => Tmkr_D0_G_negedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_G_noedge_negedge,
          SetupLow                => tsetup_D0_G_noedge_negedge,
          HoldHigh                => thold_D0_G_noedge_negedge,
          HoldLow                 => thold_D0_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( S1_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_G_negedge,
          TimingData              => Tmkr_D1_G_negedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_G_noedge_negedge,
          SetupLow                => tsetup_D1_G_noedge_negedge,
          HoldHigh                => thold_D1_G_noedge_negedge,
          HoldLow                 => thold_D1_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( S1_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_G_negedge,
          TimingData              => Tmkr_D2_G_negedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_G_noedge_negedge,
          SetupLow                => tsetup_D2_G_noedge_negedge,
          HoldHigh                => thold_D2_G_noedge_negedge,
          HoldLow                 => thold_D2_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( NOT S1_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_G_negedge,
          TimingData              => Tmkr_D3_G_negedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_G_noedge_negedge,
          SetupLow                => tsetup_D3_G_noedge_negedge,
          HoldHigh                => thold_D3_G_noedge_negedge,
          HoldLow                 => thold_D3_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( NOT S1_ipd ) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_G_negedge,
          TimingData              => Tmkr_S0_G_negedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_G_noedge_negedge,
          SetupLow                => tsetup_S0_G_noedge_negedge,
          HoldHigh                => thold_S0_G_noedge_negedge,
          HoldLow                 => thold_S0_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S1_G_negedge,
          TimingData              => Tmkr_S1_G_negedge,
          TestSignal              => S1_ipd,
          TestSignalName          => "S1",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S1_G_noedge_negedge,
          SetupLow                => tsetup_S1_G_noedge_negedge,
          HoldHigh                => thold_S1_G_noedge_negedge,
          HoldLow                 => thold_S1_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM3",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_G_negedge or Tviol_D2_G_negedge or Tviol_D3_G_negedge or Tviol_S0_G_negedge or Tviol_S1_G_negedge or Tviol_D1_G_negedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM3_Q_tab,
        DataIn => (
               D3_ipd, D2_ipd, D1_ipd, D0_ipd, S1_ipd, S0_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D0_ipd'last_event, tpd_D0_Q, TRUE),
                 1 => (D1_ipd'last_event, tpd_D1_Q, TRUE),
                 2 => (D2_ipd'last_event, tpd_D2_Q, TRUE),
                 3 => (D3_ipd'last_event, tpd_D3_Q, TRUE),
                 4 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 5 => (S1_ipd'last_event, tpd_S1_Q, TRUE),
                 6 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM3_VITAL of DLM3 is
   for VITAL_ACT
   end for;
end CFG_DLM3_VITAL;


----- CELL DLM3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S1_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S1_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM3A : entity is TRUE;
end DLM3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S1_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D0_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S1_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S1_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 6);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM3A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  L,  x,  x,  x,  L ),
    ( L,  L,  L,  x,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  L,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  H,  H,  x,  x,  x,  H ),
    ( L,  H,  H,  x,  x,  H,  x,  x,  H ),
    ( L,  H,  x,  H,  x,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  x,  L,  x,  L,  x,  L ),
    ( L,  x,  L,  x,  x,  H,  L,  x,  L ),
    ( L,  x,  H,  x,  H,  x,  L,  x,  H ),
    ( L,  x,  H,  x,  x,  H,  L,  x,  H ),
    ( L,  x,  x,  L,  L,  L,  x,  x,  L ),
    ( L,  x,  x,  L,  x,  L,  H,  x,  L ),
    ( L,  x,  x,  H,  H,  L,  x,  x,  H ),
    ( L,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( L,  x,  x,  x,  L,  L,  L,  x,  L ),
    ( L,  x,  x,  x,  H,  L,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_G_posedge,
          TimingData              => Tmkr_D0_G_posedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_G_noedge_posedge,
          SetupLow                => tsetup_D0_G_noedge_posedge,
          HoldHigh                => thold_D0_G_noedge_posedge,
          HoldLow                 => thold_D0_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( S1_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_G_posedge,
          TimingData              => Tmkr_D1_G_posedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_G_noedge_posedge,
          SetupLow                => tsetup_D1_G_noedge_posedge,
          HoldHigh                => thold_D1_G_noedge_posedge,
          HoldLow                 => thold_D1_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( S1_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_G_posedge,
          TimingData              => Tmkr_D2_G_posedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_G_noedge_posedge,
          SetupLow                => tsetup_D2_G_noedge_posedge,
          HoldHigh                => thold_D2_G_noedge_posedge,
          HoldLow                 => thold_D2_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( NOT S1_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_G_posedge,
          TimingData              => Tmkr_D3_G_posedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_G_noedge_posedge,
          SetupLow                => tsetup_D3_G_noedge_posedge,
          HoldHigh                => thold_D3_G_noedge_posedge,
          HoldLow                 => thold_D3_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( NOT S1_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_G_posedge,
          TimingData              => Tmkr_S0_G_posedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_G_noedge_posedge,
          SetupLow                => tsetup_S0_G_noedge_posedge,
          HoldHigh                => thold_S0_G_noedge_posedge,
          HoldLow                 => thold_S0_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S1_G_posedge,
          TimingData              => Tmkr_S1_G_posedge,
          TestSignal              => S1_ipd,
          TestSignalName          => "S1",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S1_G_noedge_posedge,
          SetupLow                => tsetup_S1_G_noedge_posedge,
          HoldHigh                => thold_S1_G_noedge_posedge,
          HoldLow                 => thold_S1_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM3A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_G_posedge or Tviol_S0_G_posedge or Tviol_S1_G_posedge or Tviol_D1_G_posedge or Tviol_D2_G_posedge or Tviol_D3_G_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM3A_Q_tab,
        DataIn => (
               G_ipd, D3_ipd, D2_ipd, D1_ipd, D0_ipd, S1_ipd, S0_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D0_ipd'last_event, tpd_D0_Q, TRUE),
                 1 => (D1_ipd'last_event, tpd_D1_Q, TRUE),
                 2 => (D2_ipd'last_event, tpd_D2_Q, TRUE),
                 3 => (D3_ipd'last_event, tpd_D3_Q, TRUE),
                 4 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 5 => (S1_ipd'last_event, tpd_S1_Q, TRUE),
                 6 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM3A_VITAL of DLM3A is
   for VITAL_ACT
   end for;
end CFG_DLM3A_VITAL;


----- CELL DLM4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S10_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S11_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      thold_S10_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S10_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_S11_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S11_G_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM4 : entity is TRUE;
end DLM4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S10_ipd, S11_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D0_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S10_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S10_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S11_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S11_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM4_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  H,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  x,  H,  x,  L ),
    ( L,  x,  L,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  x,  x,  x,  H,  x,  H,  H,  x,  L ),
    ( L,  x,  x,  x,  x,  H,  H,  H,  x,  L ),
    ( H,  H,  H,  H,  x,  x,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  H,  x,  x,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  H,  x,  H,  x,  H ),
    ( H,  x,  H,  x,  x,  x,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  H,  x,  H,  H,  x,  H ),
    ( H,  x,  x,  x,  x,  H,  H,  H,  x,  H ),
    ( x,  L,  x,  L,  x,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  H,  x,  L,  H,  x,  L ),
    ( x,  L,  x,  x,  x,  H,  L,  H,  x,  L ),
    ( x,  H,  x,  H,  x,  x,  L,  H,  x,  H ),
    ( x,  H,  x,  x,  H,  x,  L,  H,  x,  H ),
    ( x,  H,  x,  x,  x,  H,  L,  H,  x,  H ),
    ( x,  x,  L,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  x,  L,  x,  L,  L,  H,  H,  x,  L ),
    ( x,  x,  H,  H,  L,  L,  x,  H,  x,  H ),
    ( x,  x,  H,  x,  L,  L,  H,  H,  x,  H ),
    ( x,  x,  x,  L,  L,  L,  L,  H,  x,  L ),
    ( x,  x,  x,  H,  L,  L,  L,  H,  x,  H ),
    ( x,  x,  x,  x,  x,  x,  x,  L,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_G_negedge,
          TimingData              => Tmkr_D0_G_negedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_G_noedge_negedge,
          SetupLow                => tsetup_D0_G_noedge_negedge,
          HoldHigh                => thold_D0_G_noedge_negedge,
          HoldLow                 => thold_D0_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_G_negedge,
          TimingData              => Tmkr_D1_G_negedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_G_noedge_negedge,
          SetupLow                => tsetup_D1_G_noedge_negedge,
          HoldHigh                => thold_D1_G_noedge_negedge,
          HoldLow                 => thold_D1_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_G_negedge,
          TimingData              => Tmkr_D2_G_negedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_G_noedge_negedge,
          SetupLow                => tsetup_D2_G_noedge_negedge,
          HoldHigh                => thold_D2_G_noedge_negedge,
          HoldLow                 => thold_D2_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_G_negedge,
          TimingData              => Tmkr_D3_G_negedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_G_noedge_negedge,
          SetupLow                => tsetup_D3_G_noedge_negedge,
          HoldHigh                => thold_D3_G_noedge_negedge,
          HoldLow                 => thold_D3_G_noedge_negedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_G_negedge,
          TimingData              => Tmkr_S0_G_negedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_G_noedge_negedge,
          SetupLow                => tsetup_S0_G_noedge_negedge,
          HoldHigh                => thold_S0_G_noedge_negedge,
          HoldLow                 => thold_S0_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S10_G_negedge,
          TimingData              => Tmkr_S10_G_negedge,
          TestSignal              => S10_ipd,
          TestSignalName          => "S10",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S10_G_noedge_negedge,
          SetupLow                => tsetup_S10_G_noedge_negedge,
          HoldHigh                => thold_S10_G_noedge_negedge,
          HoldLow                 => thold_S10_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S11_G_negedge,
          TimingData              => Tmkr_S11_G_negedge,
          TestSignal              => S11_ipd,
          TestSignalName          => "S11",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S11_G_noedge_negedge,
          SetupLow                => tsetup_S11_G_noedge_negedge,
          HoldHigh                => thold_S11_G_noedge_negedge,
          HoldLow                 => thold_S11_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM4",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_G_negedge or Tviol_D2_G_negedge or Tviol_D3_G_negedge or Tviol_S0_G_negedge or Tviol_D1_G_negedge or Tviol_S10_G_negedge or Pviol_G or Tviol_S11_G_negedge;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM4_Q_tab,
        DataIn => (
               D3_ipd, D2_ipd, D1_ipd, D0_ipd, S11_ipd, S10_ipd, S0_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D0_ipd'last_event, tpd_D0_Q, TRUE),
                 1 => (D1_ipd'last_event, tpd_D1_Q, TRUE),
                 2 => (D2_ipd'last_event, tpd_D2_Q, TRUE),
                 3 => (D3_ipd'last_event, tpd_D3_Q, TRUE),
                 4 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 5 => (S10_ipd'last_event, tpd_S10_Q, TRUE),
                 6 => (S11_ipd'last_event, tpd_S11_Q, TRUE),
                 7 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM4_VITAL of DLM4 is
   for VITAL_ACT
   end for;
end CFG_DLM4_VITAL;


----- CELL DLM4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLM4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D1_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D2_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_D3_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S0_Q                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S10_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_S11_Q                      :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      thold_D0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D1_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D1_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D2_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D2_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_D3_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_D3_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S0_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S0_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      thold_S10_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S10_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_S11_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_S11_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D1                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D2                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D3                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S0                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S10                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_S11                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_G                         :	VitalDelayType01 := (1.000 ns, 1.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S10                            :	in    STD_ULOGIC;
      S11                            :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLM4A : entity is TRUE;
end DLM4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLM4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S10_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S11_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S10_ipd, S10, tipd_S10);
   VitalWireDelay (S11_ipd, S11, tipd_S11);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S10_ipd, S11_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D0_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D0_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D1_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D1_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D2_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D2_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_D3_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D3_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S0_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S0_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S10_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S10_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S11_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S11_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 7);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLM4A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  L,  x,  x,  x,  x,  L ),
    ( L,  L,  L,  x,  x,  H,  x,  x,  x,  L ),
    ( L,  L,  L,  x,  x,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  L,  x,  x,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  H,  x,  H,  x,  L ),
    ( L,  L,  x,  x,  x,  x,  H,  H,  x,  L ),
    ( L,  H,  H,  H,  H,  x,  x,  x,  x,  H ),
    ( L,  H,  H,  x,  x,  H,  x,  x,  x,  H ),
    ( L,  H,  H,  x,  x,  x,  H,  x,  x,  H ),
    ( L,  H,  x,  H,  x,  x,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  H,  x,  H,  x,  H ),
    ( L,  H,  x,  x,  x,  x,  H,  H,  x,  H ),
    ( L,  x,  L,  x,  L,  x,  x,  L,  x,  L ),
    ( L,  x,  L,  x,  x,  H,  x,  L,  x,  L ),
    ( L,  x,  L,  x,  x,  x,  H,  L,  x,  L ),
    ( L,  x,  H,  x,  H,  x,  x,  L,  x,  H ),
    ( L,  x,  H,  x,  x,  H,  x,  L,  x,  H ),
    ( L,  x,  H,  x,  x,  x,  H,  L,  x,  H ),
    ( L,  x,  x,  L,  L,  L,  L,  x,  x,  L ),
    ( L,  x,  x,  L,  x,  L,  L,  H,  x,  L ),
    ( L,  x,  x,  H,  H,  L,  L,  x,  x,  H ),
    ( L,  x,  x,  H,  x,  L,  L,  H,  x,  H ),
    ( L,  x,  x,  x,  L,  L,  L,  L,  x,  L ),
    ( L,  x,  x,  x,  H,  L,  L,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  x,  x,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D0_G_posedge,
          TimingData              => Tmkr_D0_G_posedge,
          TestSignal              => D0_ipd,
          TestSignalName          => "D0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D0_G_noedge_posedge,
          SetupLow                => tsetup_D0_G_noedge_posedge,
          HoldHigh                => thold_D0_G_noedge_posedge,
          HoldLow                 => thold_D0_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D1_G_posedge,
          TimingData              => Tmkr_D1_G_posedge,
          TestSignal              => D1_ipd,
          TestSignalName          => "D1",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D1_G_noedge_posedge,
          SetupLow                => tsetup_D1_G_noedge_posedge,
          HoldHigh                => thold_D1_G_noedge_posedge,
          HoldLow                 => thold_D1_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( S11_ipd OR S10_ipd )) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D2_G_posedge,
          TimingData              => Tmkr_D2_G_posedge,
          TestSignal              => D2_ipd,
          TestSignalName          => "D2",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D2_G_noedge_posedge,
          SetupLow                => tsetup_D2_G_noedge_posedge,
          HoldHigh                => thold_D2_G_noedge_posedge,
          HoldLow                 => thold_D2_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( S0_ipd ) OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_D3_G_posedge,
          TimingData              => Tmkr_D3_G_posedge,
          TestSignal              => D3_ipd,
          TestSignalName          => "D3",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D3_G_noedge_posedge,
          SetupLow                => tsetup_D3_G_noedge_posedge,
          HoldHigh                => thold_D3_G_noedge_posedge,
          HoldLow                 => thold_D3_G_noedge_posedge,
          CheckEnabled            => 
              TO_X01( ( NOT S0_ipd ) OR ( NOT ( S11_ipd OR S10_ipd ))) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S0_G_posedge,
          TimingData              => Tmkr_S0_G_posedge,
          TestSignal              => S0_ipd,
          TestSignalName          => "S0",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S0_G_noedge_posedge,
          SetupLow                => tsetup_S0_G_noedge_posedge,
          HoldHigh                => thold_S0_G_noedge_posedge,
          HoldLow                 => thold_S0_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S10_G_posedge,
          TimingData              => Tmkr_S10_G_posedge,
          TestSignal              => S10_ipd,
          TestSignalName          => "S10",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S10_G_noedge_posedge,
          SetupLow                => tsetup_S10_G_noedge_posedge,
          HoldHigh                => thold_S10_G_noedge_posedge,
          HoldLow                 => thold_S10_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S11_G_posedge,
          TimingData              => Tmkr_S11_G_posedge,
          TestSignal              => S11_ipd,
          TestSignalName          => "S11",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S11_G_noedge_posedge,
          SetupLow                => tsetup_S11_G_noedge_posedge,
          HoldHigh                => thold_S11_G_noedge_posedge,
          HoldLow                 => thold_S11_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLM4A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D0_G_posedge or Tviol_S0_G_posedge or Tviol_D1_G_posedge or Tviol_D2_G_posedge or Tviol_D3_G_posedge or Tviol_S10_G_posedge or Tviol_S11_G_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLM4A_Q_tab,
        DataIn => (
               G_ipd, D3_ipd, D2_ipd, D1_ipd, D0_ipd, S11_ipd, S10_ipd, S0_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D0_ipd'last_event, tpd_D0_Q, TRUE),
                 1 => (D1_ipd'last_event, tpd_D1_Q, TRUE),
                 2 => (D2_ipd'last_event, tpd_D2_Q, TRUE),
                 3 => (D3_ipd'last_event, tpd_D3_Q, TRUE),
                 4 => (S0_ipd'last_event, tpd_S0_Q, TRUE),
                 5 => (S10_ipd'last_event, tpd_S10_Q, TRUE),
                 6 => (S11_ipd'last_event, tpd_S11_Q, TRUE),
                 7 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLM4A_VITAL of DLM4A is
   for VITAL_ACT
   end for;
end CFG_DLM4A_VITAL;


----- CELL DLMA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLMA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLMA : entity is TRUE;
end DLMA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLMA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_A_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 3);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLMA_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  x,  L ),
    ( L,  L,  x,  H,  x,  L ),
    ( L,  H,  H,  x,  x,  H ),
    ( L,  H,  x,  H,  x,  H ),
    ( L,  x,  L,  L,  x,  L ),
    ( L,  x,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_G_posedge,
          TimingData              => Tmkr_A_G_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_G_noedge_posedge,
          SetupLow                => tsetup_A_G_noedge_posedge,
          HoldHigh                => thold_A_G_noedge_posedge,
          HoldLow                 => thold_A_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( ( S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_G_posedge,
          TimingData              => Tmkr_B_G_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_G_noedge_posedge,
          SetupLow                => tsetup_B_G_noedge_posedge,
          HoldHigh                => thold_B_G_noedge_posedge,
          HoldLow                 => thold_B_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01( (NOT S_ipd ) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_G_posedge,
          TimingData              => Tmkr_S_G_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_G_noedge_posedge,
          SetupLow                => tsetup_S_G_noedge_posedge,
          HoldHigh                => thold_S_G_noedge_posedge,
          HoldLow                 => thold_S_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLMA",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_G_posedge or Tviol_B_G_posedge or Tviol_S_G_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLMA_Q_tab,
        DataIn => (
               G_ipd, B_ipd, A_ipd, S_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE),
                 3 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLMA_VITAL of DLMA is
   for VITAL_ACT
   end for;
end CFG_DLMA_VITAL;


----- CELL DLME1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLME1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_A_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_A_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_A_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_A_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_B_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_B_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_B_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_B_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_S_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      thold_S_E_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_S_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tsetup_S_E_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_E_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLME1A : entity is TRUE;
end DLME1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLME1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd, E_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_A_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_A_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_A_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_B_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_B_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_S_E_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_S_E_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_E	: STD_ULOGIC := '0';
   VARIABLE PInfo_E	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLME1A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  L,  x,  x,  L ),
    ( L,  L,  L,  x,  H,  x,  L ),
    ( L,  L,  H,  H,  x,  x,  H ),
    ( L,  L,  H,  x,  H,  x,  H ),
    ( L,  L,  x,  L,  L,  x,  L ),
    ( L,  L,  x,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  x,  S ),
    ( x,  H,  x,  x,  x,  x,  S ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_A_G_posedge,
          TimingData              => Tmkr_A_G_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_G_noedge_posedge,
          SetupLow                => tsetup_A_G_noedge_posedge,
          HoldHigh                => thold_A_G_noedge_posedge,
          HoldLow                 => thold_A_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(E_ipd OR S_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_A_E_posedge,
          TimingData              => Tmkr_A_E_posedge,
          TestSignal              => A_ipd,
          TestSignalName          => "A",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_A_E_noedge_posedge,
          SetupLow                => tsetup_A_E_noedge_posedge,
          HoldHigh                => thold_A_E_noedge_posedge,
          HoldLow                 => thold_A_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(S_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_G_posedge,
          TimingData              => Tmkr_B_G_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_G_noedge_posedge,
          SetupLow                => tsetup_B_G_noedge_posedge,
          HoldHigh                => thold_B_G_noedge_posedge,
          HoldLow                 => thold_B_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(E_ipd OR (NOT S_ipd)) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_B_E_posedge,
          TimingData              => Tmkr_B_E_posedge,
          TestSignal              => B_ipd,
          TestSignalName          => "B",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_B_E_noedge_posedge,
          SetupLow                => tsetup_B_E_noedge_posedge,
          HoldHigh                => thold_B_E_noedge_posedge,
          HoldLow                 => thold_B_E_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(NOT S_ipd) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_G_posedge,
          TimingData              => Tmkr_S_G_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_G_noedge_posedge,
          SetupLow                => tsetup_S_G_noedge_posedge,
          HoldHigh                => thold_S_G_noedge_posedge,
          HoldLow                 => thold_S_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_S_E_posedge,
          TimingData              => Tmkr_S_E_posedge,
          TestSignal              => S_ipd,
          TestSignalName          => "S",
          TestDelay               => 0 ns,
          RefSignal               => E_ipd,
          RefSignalName          => "E",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_S_E_noedge_posedge,
          SetupLow                => tsetup_S_E_noedge_posedge,
          HoldHigh                => thold_S_E_noedge_posedge,
          HoldLow                 => thold_S_E_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_E,
          PeriodData              => PInfo_E,
          TestSignal              => E_ipd,
          TestSignalName          => "E",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_E_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLME1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_A_G_posedge or Pviol_E or Tviol_A_E_posedge or Tviol_B_G_posedge or Tviol_B_E_posedge or Tviol_S_G_posedge or Tviol_S_E_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLME1A_Q_tab,
        DataIn => (
               G_ipd, E_ipd, B_ipd, A_ipd, S_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Q, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Q, TRUE),
                 2 => (S_ipd'last_event, tpd_S_Q, TRUE),
                 3 => (E_ipd'last_event, tpd_E_Q, TRUE),
                 4 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLME1A_VITAL of DLME1A is
   for VITAL_ACT
   end for;
end CFG_DLME1A_VITAL;


----- CELL DLP1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLP1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLP1 : entity is TRUE;
end DLP1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLP1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLP1_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( H,  x,  H,  x,  H ),
    ( x,  L,  L,  x,  S ),
    ( x,  H,  x,  x,  H ),
    ( x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_negedge,
          TimingData              => Tmkr_PRE_G_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_negedge_negedge,
          Removal                 => thold_PRE_G_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLP1",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLP1_Q_tab,
        DataIn => (
               D_ipd, PRE_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLP1_VITAL of DLP1 is
   for VITAL_ACT
   end for;
end CFG_DLP1_VITAL;


----- CELL DLP1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLP1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_negedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_PRE_posedge                :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLP1A : entity is TRUE;
end DLP1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLP1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLP1A_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  L ),
    ( L,  H,  x,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  x,  H,  x,  H ),
    ( x,  x,  U,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_posedge,
          TimingData              => Tmkr_PRE_G_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_negedge_posedge,
          Removal                 => thold_PRE_G_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01(PRE_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/DLP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_PRE_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLP1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLP1A_Q_tab,
        DataIn => (
               G_ipd, D_ipd, PRE_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLP1A_VITAL of DLP1A is
   for VITAL_ACT
   end for;
end CFG_DLP1A_VITAL;


----- CELL DLP1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLP1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLP1B : entity is TRUE;
end DLP1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLP1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLP1B_Q_tab : VitalStateTableType := (
    ( L,  H,  H,  x,  L ),
    ( H,  x,  H,  x,  H ),
    ( x,  L,  x,  x,  H ),
    ( x,  H,  L,  x,  S ),
    ( x,  U,  x,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_negedge,
          TimingData              => Tmkr_PRE_G_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_posedge_negedge,
          Removal                 => thold_PRE_G_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLP1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLP1B_Q_tab,
        DataIn => (
               D_ipd, PRE_ipd, G_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLP1B_VITAL of DLP1B is
   for VITAL_ACT
   end for;
end CFG_DLP1B_VITAL;


----- CELL DLP1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLP1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLP1C : entity is TRUE;
end DLP1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLP1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLP1C_Q_tab : VitalStateTableType := (
    ( L,  L,  H,  x,  L ),
    ( L,  H,  x,  x,  H ),
    ( H,  x,  H,  x,  S ),
    ( x,  x,  L,  x,  H ),
    ( x,  x,  U,  H,  H ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_posedge,
          TimingData              => Tmkr_PRE_G_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_posedge_posedge,
          Removal                 => thold_PRE_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLP1C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DLP1C_Q_tab,
        DataIn => (
               G_ipd, D_ipd, PRE_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLP1C_VITAL of DLP1C is
   for VITAL_ACT
   end for;
end CFG_DLP1C_VITAL;


----- CELL DLP1D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLP1D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_negedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_negedge              :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLP1D : entity is TRUE;
end DLP1D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLP1D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLP1D_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  L,  H,  x,  H ),
    ( H,  x,  L,  x,  S ),
    ( x,  H,  H,  x,  L ),
    ( U,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_negedge,
          TimingData              => Tmkr_PRE_G_negedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_posedge_negedge,
          Removal                 => thold_PRE_G_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/DLP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_negedge,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLP1D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Tviol_PRE_G_negedge or Pviol_PRE or Pviol_G;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DLP1D_QN_tab,
        DataIn => (
               PRE_ipd, D_ipd, G_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLP1D_VITAL of DLP1D is
   for VITAL_ACT
   end for;
end CFG_DLP1D_VITAL;


----- CELL DLP1E -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DLP1E is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_QN                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_PRE_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_posedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_posedge                     :	VitalDelayType := 0.000 ns;
      thold_PRE_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      trecovery_PRE_G_posedge_posedge                :	VitalDelayType := 0.000 ns;
      tperiod_G_posedge              :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tpw_PRE_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_PRE                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PRE                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DLP1E : entity is TRUE;
end DLP1E;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of DLP1E is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL PRE_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (PRE_ipd, PRE, tipd_PRE);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd, PRE_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_PRE_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PRE_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_PRE	: STD_ULOGIC := '0';
   VARIABLE PInfo_PRE	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DLP1E_QN_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  L ),
    ( H,  L,  L,  x,  H ),
    ( H,  H,  x,  x,  S ),
    ( x,  L,  H,  x,  L ),
    ( U,  x,  x,  L,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_posedge,
          TimingData              => Tmkr_D_G_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_posedge,
          SetupLow                => tsetup_D_G_noedge_posedge,
          HoldHigh                => thold_D_G_noedge_posedge,
          HoldLow                 => thold_D_G_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_PRE_G_posedge,
          TimingData              => Tmkr_PRE_G_posedge,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          Recovery                => trecovery_PRE_G_posedge_posedge,
          Removal                 => thold_PRE_G_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/DLP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => tperiod_G_posedge,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TO_X01((NOT PRE_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/DLP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_PRE,
          PeriodData              => PInfo_PRE,
          TestSignal              => PRE_ipd,
          TestSignalName          => "PRE",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_PRE_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/DLP1E",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_posedge or Tviol_PRE_G_posedge or Pviol_PRE or Pviol_G;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DLP1E_QN_tab,
        DataIn => (
               PRE_ipd, G_ipd, D_ipd));
      QN_zd := Violation XOR QN_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_QN, TRUE),
                 1 => (G_ipd'last_event, tpd_G_QN, TRUE),
                 2 => (PRE_ipd'last_event, tpd_PRE_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DLP1E_VITAL of DLP1E is
   for VITAL_ACT
   end for;
end CFG_DLP1E_VITAL;


----- CELL DXAND7 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DXAND7 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_F_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_F                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      F                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DXAND7 : entity is TRUE;
end DXAND7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DXAND7 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL F_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (F_ipd, F, tipd_F);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd, F_ipd, G_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (B_ipd) AND (A_ipd) AND (C_ipd) AND (D_ipd) AND (E_ipd) AND (F_ipd)
         AND (G_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 1 => (F_ipd'last_event, tpd_F_Y, TRUE),
                 2 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 5 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 6 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DXAND7_VITAL of DXAND7 is
   for VITAL_ACT
   end for;
end CFG_DXAND7_VITAL;


----- CELL DXAX7 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DXAX7 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_H_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_F_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_F                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_H                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      F                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      H                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DXAX7 : entity is TRUE;
end DXAX7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DXAX7 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL F_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';
   SIGNAL H_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (F_ipd, F, tipd_F);
   VitalWireDelay (G_ipd, G, tipd_G);
   VitalWireDelay (H_ipd, H, tipd_H);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd, F_ipd, G_ipd, H_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (H_ipd) XOR ((B_ipd) AND (A_ipd) AND (C_ipd) AND (D_ipd) AND (E_ipd)
         AND (F_ipd) AND (G_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (H_ipd'last_event, tpd_H_Y, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 2 => (F_ipd'last_event, tpd_F_Y, TRUE),
                 3 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 4 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 5 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 6 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 7 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DXAX7_VITAL of DXAX7 is
   for VITAL_ACT
   end for;
end CFG_DXAX7_VITAL;


----- CELL DXNAND7 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity DXNAND7 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_F_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_F                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      F                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of DXNAND7 : entity is TRUE;
end DXNAND7;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of DXNAND7 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL F_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (F_ipd, F, tipd_F);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd, F_ipd, G_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT ((B_ipd) AND (A_ipd) AND (C_ipd) AND (D_ipd) AND (E_ipd) AND
         (F_ipd) AND (G_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 1 => (F_ipd'last_event, tpd_F_Y, TRUE),
                 2 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 5 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 6 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_DXNAND7_VITAL of DXNAND7 is
   for VITAL_ACT
   end for;
end CFG_DXNAND7_VITAL;


----- CELL FA1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity FA1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CI_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CI_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CI                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CI                             :	in    STD_ULOGIC;
      S                              :	out   STD_ULOGIC;
      CO                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of FA1A : entity is TRUE;
end FA1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of FA1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CI_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (CI_ipd, CI, tipd_CI);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, CI_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS S_zd : STD_LOGIC is Results(1);
   ALIAS CO_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE S_GlitchData	: VitalGlitchDataType;
   VARIABLE CO_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      S_zd :=
       (((NOT A_ipd)) AND ((((NOT B_ipd)) AND (A_ipd)) OR (((NOT B_ipd)) AND
         (CI_ipd) AND ((NOT A_ipd))) OR ((CI_ipd) AND (B_ipd) AND (A_ipd)))
         AND (CI_ipd)) OR (((NOT A_ipd)) AND (B_ipd) AND ((NOT CI_ipd))) OR
         ((A_ipd) AND ((((NOT B_ipd)) AND (A_ipd)) OR (((NOT B_ipd)) AND
         (CI_ipd) AND ((NOT A_ipd))) OR ((CI_ipd) AND (B_ipd) AND (A_ipd)))
         AND ((NOT CI_ipd))) OR ((A_ipd) AND (B_ipd) AND (CI_ipd));
      CO_zd :=
       (((NOT B_ipd)) AND (A_ipd)) OR (((NOT B_ipd)) AND (CI_ipd)) OR 
       ((CI_ipd) AND (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (CI_ipd'last_event, tpd_CI_S, TRUE),
                 1 => (B_ipd'last_event, tpd_B_S, TRUE),
                 2 => (A_ipd'last_event, tpd_A_S, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (CI_ipd'last_event, tpd_CI_CO, TRUE),
                 1 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 2 => (A_ipd'last_event, tpd_A_CO, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_FA1A_VITAL of FA1A is
   for VITAL_ACT
   end for;
end CFG_FA1A_VITAL;


----- CELL FA1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity FA1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CI_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CI_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CI                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CI                             :	in    STD_ULOGIC;
      S                              :	out   STD_ULOGIC;
      CO                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of FA1B : entity is TRUE;
end FA1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of FA1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CI_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (CI_ipd, CI, tipd_CI);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, CI_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS S_zd : STD_LOGIC is Results(1);
   ALIAS CO_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE S_GlitchData	: VitalGlitchDataType;
   VARIABLE CO_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      S_zd :=
       ((((((CI_ipd) AND ((NOT B_ipd)) AND (A_ipd)) OR ((((CI_ipd) AND
         (B_ipd)) OR ((NOT B_ipd))) AND ((NOT A_ipd)))) AND (CI_ipd)) OR
         ((B_ipd) AND ((NOT CI_ipd)))) AND (A_ipd)) OR ((((B_ipd) AND
         (CI_ipd)) OR ((((CI_ipd) AND ((NOT B_ipd)) AND (A_ipd)) OR
         ((((CI_ipd) AND (B_ipd)) OR ((NOT B_ipd))) AND ((NOT A_ipd)))) AND
         ((NOT CI_ipd)))) AND ((NOT A_ipd)));
      CO_zd :=
       ((CI_ipd) AND ((NOT B_ipd))) OR ((CI_ipd) AND ((NOT A_ipd)))
         OR (((NOT B_ipd)) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (CI_ipd'last_event, tpd_CI_S, TRUE),
                 1 => (B_ipd'last_event, tpd_B_S, TRUE),
                 2 => (A_ipd'last_event, tpd_A_S, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (CI_ipd'last_event, tpd_CI_CO, TRUE),
                 1 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 2 => (A_ipd'last_event, tpd_A_CO, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_FA1B_VITAL of FA1B is
   for VITAL_ACT
   end for;
end CFG_FA1B_VITAL;


----- CELL FA2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity FA2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CI_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_S                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CI_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A1_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A0_CO                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_A1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CI                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A0                             :	in    STD_ULOGIC;
      A1                             :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CI                             :	in    STD_ULOGIC;
      S                              :	out   STD_ULOGIC;
      CO                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of FA2A : entity is TRUE;
end FA2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of FA2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL A1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CI_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A0_ipd, A0, tipd_A0);
   VitalWireDelay (A1_ipd, A1, tipd_A1);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (CI_ipd, CI, tipd_CI);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A0_ipd, A1_ipd, B_ipd, CI_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS S_zd : STD_LOGIC is Results(1);
   ALIAS CO_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE S_GlitchData	: VitalGlitchDataType;
   VARIABLE CO_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      S_zd :=
       (((NOT ((A1_ipd) OR (A0_ipd)))) AND ((((A1_ipd) OR (A0_ipd)) AND
         ((NOT B_ipd))) OR (((NOT B_ipd)) AND (CI_ipd) AND ((NOT ((A1_ipd) OR
         (A0_ipd))))) OR ((CI_ipd) AND (B_ipd) AND ((A1_ipd) OR (A0_ipd))))
         AND (CI_ipd)) OR (((NOT ((A1_ipd) OR (A0_ipd)))) AND (B_ipd) AND
         ((NOT CI_ipd))) OR (((A1_ipd) OR (A0_ipd)) AND ((((A1_ipd) OR
         (A0_ipd)) AND ((NOT B_ipd))) OR (((NOT B_ipd)) AND (CI_ipd) AND
         ((NOT ((A1_ipd) OR (A0_ipd))))) OR ((CI_ipd) AND (B_ipd) AND
         ((A1_ipd) OR (A0_ipd)))) AND ((NOT CI_ipd))) OR (((A1_ipd) OR
         (A0_ipd)) AND (B_ipd) AND (CI_ipd));
      --CO_zd :=
      -- (((A1_ipd) OR (A0_ipd)) AND ((NOT B_ipd))) OR (((NOT B_ipd)) AND
      --   (CI_ipd) AND ((NOT ((A1_ipd) OR (A0_ipd))))) OR ((CI_ipd) AND
      --   (B_ipd) AND ((A1_ipd) OR (A0_ipd)));
      CO_zd := 
        (((A1_ipd) AND (NOT B_ipd)) OR ((A0_ipd) AND (NOT B_ipd)) OR
         ((A0_ipd) AND (CI_ipd)) OR ((A1_ipd) AND (CI_ipd)) OR
         ((NOT B_ipd) AND (CI_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (CI_ipd'last_event, tpd_CI_S, TRUE),
                 1 => (B_ipd'last_event, tpd_B_S, TRUE),
                 2 => (A1_ipd'last_event, tpd_A1_S, TRUE),
                 3 => (A0_ipd'last_event, tpd_A0_S, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (CI_ipd'last_event, tpd_CI_CO, TRUE),
                 1 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 2 => (A1_ipd'last_event, tpd_A1_CO, TRUE),
                 3 => (A0_ipd'last_event, tpd_A0_CO, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_FA2A_VITAL of FA2A is
   for VITAL_ACT
   end for;
end CFG_FA2A_VITAL;


----- CELL GAND2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GAND2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of GAND2 : entity is TRUE;
end GAND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of GAND2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, G_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (G_ipd) AND (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_GAND2_VITAL of GAND2 is
   for VITAL_ACT
   end for;
end CFG_GAND2_VITAL;


----- CELL GMX4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GMX4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of GMX4 : entity is TRUE;
end GMX4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of GMX4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, G_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := VitalMUX
                 (data => (D3_ipd, D1_ipd, D2_ipd, D0_ipd),
                  dselect => (S0_ipd, G_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 1 => (S0_ipd'last_event, tpd_S0_Y, TRUE),
                 2 => (D3_ipd'last_event, tpd_D3_Y, TRUE),
                 3 => (D2_ipd'last_event, tpd_D2_Y, TRUE),
                 4 => (D1_ipd'last_event, tpd_D1_Y, TRUE),
                 5 => (D0_ipd'last_event, tpd_D0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_GMX4_VITAL of GMX4 is
   for VITAL_ACT
   end for;
end CFG_GMX4_VITAL;


----- CELL GNAND2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GNAND2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of GNAND2 : entity is TRUE;
end GNAND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of GNAND2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, G_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((G_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_GNAND2_VITAL of GNAND2 is
   for VITAL_ACT
   end for;
end CFG_GNAND2_VITAL;


----- CELL GND -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GND is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True);

   port(
      Y                              :	out   STD_ULOGIC := '0');
attribute VITAL_LEVEL0 of GND : entity is TRUE;
end GND;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of GND is
   attribute VITAL_LEVEL0 of VITAL_ACT : architecture is TRUE;


begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   --  empty
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   Y <= '0';



end VITAL_ACT;

configuration CFG_GND_VITAL of GND is
   for VITAL_ACT
   end for;
end CFG_GND_VITAL;



----- CELL GNOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GNOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of GNOR2 : entity is TRUE;
end GNOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of GNOR2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, G_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((G_ipd) OR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_GNOR2_VITAL of GNOR2 is
   for VITAL_ACT
   end for;
end CFG_GNOR2_VITAL;


----- CELL GOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of GOR2 : entity is TRUE;
end GOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of GOR2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, G_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (G_ipd) OR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_GOR2_VITAL of GOR2 is
   for VITAL_ACT
   end for;
end CFG_GOR2_VITAL;


----- CELL GXOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity GXOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_G_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of GXOR2 : entity is TRUE;
end GXOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of GXOR2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, G_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (G_ipd) XOR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (G_ipd'last_event, tpd_G_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_GXOR2_VITAL of GXOR2 is
   for VITAL_ACT
   end for;
end CFG_GXOR2_VITAL;


----- CELL HA1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity HA1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of HA1 : entity is TRUE;
end HA1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of HA1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS CO_zd : STD_LOGIC is Results(1);
   ALIAS S_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE CO_GlitchData	: VitalGlitchDataType;
   VARIABLE S_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      CO_zd := (B_ipd) AND (A_ipd);
      S_zd := (B_ipd) XOR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 1 => (A_ipd'last_event, tpd_A_CO, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_S, TRUE),
                 1 => (A_ipd'last_event, tpd_A_S, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_HA1_VITAL of HA1 is
   for VITAL_ACT
   end for;
end CFG_HA1_VITAL;


----- CELL HA1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity HA1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of HA1A : entity is TRUE;
end HA1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of HA1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS CO_zd : STD_LOGIC is Results(1);
   ALIAS S_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE CO_GlitchData	: VitalGlitchDataType;
   VARIABLE S_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      CO_zd := (B_ipd) AND ((NOT A_ipd));
      S_zd := (NOT ((B_ipd) XOR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 1 => (A_ipd'last_event, tpd_A_CO, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_S, TRUE),
                 1 => (A_ipd'last_event, tpd_A_S, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_HA1A_VITAL of HA1A is
   for VITAL_ACT
   end for;
end CFG_HA1A_VITAL;


----- CELL HA1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity HA1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of HA1B : entity is TRUE;
end HA1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of HA1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS CO_zd : STD_LOGIC is Results(1);
   ALIAS S_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE CO_GlitchData	: VitalGlitchDataType;
   VARIABLE S_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      CO_zd := (NOT ((B_ipd) AND (A_ipd)));
      S_zd := (NOT ((B_ipd) XOR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 1 => (A_ipd'last_event, tpd_A_CO, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_S, TRUE),
                 1 => (A_ipd'last_event, tpd_A_S, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_HA1B_VITAL of HA1B is
   for VITAL_ACT
   end for;
end CFG_HA1B_VITAL;


----- CELL HA1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity HA1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_CO                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_S                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      CO                             :	out   STD_ULOGIC;
      S                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of HA1C : entity is TRUE;
end HA1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of HA1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 2) := (others => 'X');
   ALIAS CO_zd : STD_LOGIC is Results(1);
   ALIAS S_zd : STD_LOGIC is Results(2);

   -- output glitch detection variables
   VARIABLE CO_GlitchData	: VitalGlitchDataType;
   VARIABLE S_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      CO_zd := (NOT ((B_ipd) AND (A_ipd)));
      S_zd := (B_ipd) XOR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => CO,
       GlitchData => CO_GlitchData,
       OutSignalName => "CO",
       OutTemp => CO_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_CO, TRUE),
                 1 => (A_ipd'last_event, tpd_A_CO, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);
      VitalPathDelay01 (
       OutSignal => S,
       GlitchData => S_GlitchData,
       OutSignalName => "S",
       OutTemp => S_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_S, TRUE),
                 1 => (A_ipd'last_event, tpd_A_S, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_HA1C_VITAL of HA1C is
   for VITAL_ACT
   end for;
end CFG_HA1C_VITAL;


----- CELL IBDL -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IBDL is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_Q                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_PAD_G_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_PAD_G_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_G_negedge                  :	VitalDelayType := 0.000 ns;
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IBDL : entity is TRUE;
end IBDL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of IBDL is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_PAD_G_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PAD_G_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_PAD_G_posedge,
          TimingData              => Tmkr_PAD_G_posedge,
          TestSignal              => PAD_ipd,
          TestSignalName          => "PAD",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_PAD_G_noedge_posedge,
          SetupLow                => tsetup_PAD_G_noedge_posedge,
          HoldHigh                => thold_PAD_G_noedge_posedge,
          HoldLow                 => thold_PAD_G_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IBDL",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_G_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/IBDL",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_PAD_G_posedge or Pviol_G;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DL1B_Q_tab,
        DataIn => (
               G_ipd, PAD_ipd));
      Q_zd := Violation XOR Q_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Q, TRUE),
                 1 => (G_ipd'last_event, tpd_G_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IBDL_VITAL of IBDL is
   for VITAL_ACT
   end for;
end CFG_IBDL_VITAL;


----- CELL INBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INBUF : entity is TRUE;
end INBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of INBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_INBUF_VITAL of INBUF is
   for VITAL_ACT
   end for;
end CFG_INBUF_VITAL;


----- CELL INV -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INV is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INV : entity is TRUE;
end INV;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of INV is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_INV_VITAL of INV is
   for VITAL_ACT
   end for;
end CFG_INV_VITAL;


----- CELL INVA -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INVA is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INVA : entity is TRUE;
end INVA;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of INVA is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_INVA_VITAL of INVA is
   for VITAL_ACT
   end for;
end CFG_INVA_VITAL;


----- CELL INVD -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity INVD is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of INVD : entity is TRUE;
end INVD;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of INVD is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_INVD_VITAL of INVD is
   for VITAL_ACT
   end for;
end CFG_INVD_VITAL;


----- CELL IR -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IR is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_PAD_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_PAD_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IR : entity is TRUE;
end IR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of IR is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_PAD_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PAD_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE PAD_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_PAD_CLK_posedge,
          TimingData              => Tmkr_PAD_CLK_posedge,
          TestSignal              => PAD_ipd,
          TestSignalName          => "PAD",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_PAD_CLK_noedge_posedge,
          SetupLow                => tsetup_PAD_CLK_noedge_posedge,
          HoldHigh                => thold_PAD_CLK_noedge_posedge,
          HoldLow                 => thold_PAD_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/IR",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_PAD_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DF1_Q_tab,
        DataIn => (
               CLK_delayed, PAD_delayed, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      PAD_delayed := PAD_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IR_VITAL of IR is
   for VITAL_ACT
   end for;
end CFG_IR_VITAL;


----- CELL IRI -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity IRI is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_QN                     :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_PAD_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      tsetup_PAD_CLK_noedge_posedge                 :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      QN                             :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of IRI : entity is TRUE;
end IRI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of IRI is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_PAD_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_PAD_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_QN : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE PAD_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS QN_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE QN_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_PAD_CLK_posedge,
          TimingData              => Tmkr_PAD_CLK_posedge,
          TestSignal              => PAD_ipd,
          TestSignalName          => "PAD",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_PAD_CLK_noedge_posedge,
          SetupLow                => tsetup_PAD_CLK_noedge_posedge,
          HoldHigh                => thold_PAD_CLK_noedge_posedge,
          HoldLow                 => thold_PAD_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/IRI",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/IRI",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_PAD_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => QN_zd,
        PreviousDataIn => PrevData_QN,
        StateTable => DF1A_QN_tab,
        DataIn => (
               CLK_delayed, PAD_delayed, CLK_ipd));
      QN_zd := Violation XOR QN_zd;
      PAD_delayed := PAD_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => QN,
       GlitchData => QN_GlitchData,
       OutSignalName => "QN",
       OutTemp => QN_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QN, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_IRI_VITAL of IRI is
   for VITAL_ACT
   end for;
end CFG_IRI_VITAL;


----- CELL JKF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKF : entity is TRUE;
end JKF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of JKF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (J_ipd, K_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_J_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_posedge,
          TimingData              => Tmkr_J_CLK_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_posedge,
          TimingData              => Tmkr_K_CLK_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKF",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_posedge or Tviol_K_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_delayed, K_delayed, J_delayed, Q_zd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_JKF_VITAL of JKF is
   for VITAL_ACT
   end for;
end CFG_JKF_VITAL;


----- CELL JKF1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKF1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKF1B : entity is TRUE;
end JKF1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of JKF1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (J_ipd, K_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_J_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_negedge,
          TimingData              => Tmkr_J_CLK_negedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_J_CLK_noedge_negedge,
          SetupLow                => tsetup_J_CLK_noedge_negedge,
          HoldHigh                => thold_J_CLK_noedge_negedge,
          HoldLow                 => thold_J_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_negedge,
          TimingData              => Tmkr_K_CLK_negedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_K_CLK_noedge_negedge,
          SetupLow                => tsetup_K_CLK_noedge_negedge,
          HoldHigh                => thold_K_CLK_noedge_negedge,
          HoldLow                 => thold_K_CLK_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_negedge or Tviol_K_CLK_negedge or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE1B_Q_tab,
        DataIn => (
               CLK_ipd, K_delayed, J_delayed, Q_zd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_JKF1B_VITAL of JKF1B is
   for VITAL_ACT
   end for;
end CFG_JKF1B_VITAL;


----- CELL JKF2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKF2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKF2A : entity is TRUE;
end JKF2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of JKF2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (J_ipd, K_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_J_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_posedge,
          TimingData              => Tmkr_J_CLK_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_posedge,
          TimingData              => Tmkr_K_CLK_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/JKF2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKF2A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_posedge or Tviol_CLR_CLK_posedge or Tviol_K_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, K_delayed, J_delayed, Q_zd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_JKF2A_VITAL of JKF2A is
   for VITAL_ACT
   end for;
end CFG_JKF2A_VITAL;


----- CELL JKF2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKF2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKF2B : entity is TRUE;
end JKF2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of JKF2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (J_ipd, K_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_J_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFE3C_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  H,  H,  x,  H,  x,  H ),
    ( H,  L,  H,  x,  H,  H,  x,  H ),
    ( H,  L,  x,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  x,  H,  x,  L ),
    ( x,  L,  L,  x,  H,  H,  x,  L ),
    ( x,  L,  x,  L,  L,  H,  x,  L ),
    ( U,  x,  x,  x,  L,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_negedge,
          TimingData              => Tmkr_J_CLK_negedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_J_CLK_noedge_negedge,
          SetupLow                => tsetup_J_CLK_noedge_negedge,
          HoldHigh                => thold_J_CLK_noedge_negedge,
          HoldLow                 => thold_J_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_negedge,
          TimingData              => Tmkr_K_CLK_negedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_K_CLK_noedge_negedge,
          SetupLow                => tsetup_K_CLK_noedge_negedge,
          HoldHigh                => thold_K_CLK_noedge_negedge,
          HoldLow                 => thold_K_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/JKF2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKF2B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_negedge or Tviol_K_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFE3C_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, K_delayed, J_delayed, Q_zd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_JKF2B_VITAL of JKF2B is
   for VITAL_ACT
   end for;
end CFG_JKF2B_VITAL;


----- CELL JKF2C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKF2C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKF2C : entity is TRUE;
end JKF2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of JKF2C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (J_ipd, K_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_J_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM3_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  x,  L ),
    ( L,  H,  H,  x,  H,  L,  x,  H ),
    ( L,  H,  x,  H,  H,  L,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  x,  L ),
    ( L,  x,  H,  L,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  x,  x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  L,  x,  U,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_posedge,
          TimingData              => Tmkr_J_CLK_posedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_J_CLK_noedge_posedge,
          SetupLow                => tsetup_J_CLK_noedge_posedge,
          HoldHigh                => thold_J_CLK_noedge_posedge,
          HoldLow                 => thold_J_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_posedge,
          TimingData              => Tmkr_K_CLK_posedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_K_CLK_noedge_posedge,
          SetupLow                => tsetup_K_CLK_noedge_posedge,
          HoldHigh                => thold_K_CLK_noedge_posedge,
          HoldLow                 => thold_K_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/JKF2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/JKF2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKF2C",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_posedge or Tviol_CLR_CLK_posedge or Tviol_K_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM3_Q_tab,
        DataIn => (
               CLK_delayed, K_delayed, J_delayed, Q_zd, CLK_ipd, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_JKF2C_VITAL of JKF2C is
   for VITAL_ACT
   end for;
end CFG_JKF2C_VITAL;


----- CELL JKF2D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity JKF2D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_J_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_J_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_K_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_K_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_negedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_J                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_K                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      J                              :	in    STD_ULOGIC;
      K                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of JKF2D : entity is TRUE;
end JKF2D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of JKF2D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL J_ipd	 : STD_ULOGIC := 'X';
   SIGNAL K_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (J_ipd, J, tipd_J);
   VitalWireDelay (K_ipd, K, tipd_K);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (J_ipd, K_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_J_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_J_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_K_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_K_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 5);
   VARIABLE J_delayed : STD_ULOGIC := 'X';
   VARIABLE K_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT DFM3_Q_tab : VitalStateTableType := (
    ( L,  L,  L,  x,  H,  x,  x,  L ),
    ( L,  L,  x,  H,  H,  x,  x,  L ),
    ( L,  H,  H,  x,  H,  L,  x,  H ),
    ( L,  H,  x,  H,  H,  L,  x,  H ),
    ( L,  x,  L,  L,  H,  x,  x,  L ),
    ( L,  x,  H,  L,  H,  L,  x,  H ),
    ( H,  x,  x,  x,  x,  L,  x,  S ),
    ( x,  x,  x,  x,  L,  L,  x,  S ),
    ( x,  x,  x,  x,  x,  H,  x,  L ),
    ( x,  x,  x,  L,  x,  U,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_J_CLK_negedge,
          TimingData              => Tmkr_J_CLK_negedge,
          TestSignal              => J_ipd,
          TestSignalName          => "J",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_J_CLK_noedge_negedge,
          SetupLow                => tsetup_J_CLK_noedge_negedge,
          HoldHigh                => thold_J_CLK_noedge_negedge,
          HoldLow                 => thold_J_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalSetupHoldCheck (
          Violation               => Tviol_K_CLK_negedge,
          TimingData              => Tmkr_K_CLK_negedge,
          TestSignal              => K_ipd,
          TestSignalName          => "K",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_K_CLK_noedge_negedge,
          SetupLow                => tsetup_K_CLK_noedge_negedge,
          HoldHigh                => thold_K_CLK_noedge_negedge,
          HoldLow                 => thold_K_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_negedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => FALSE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/JKF2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01(CLR_ipd ) /= '1',
          HeaderMsg               => InstancePath &"/JKF2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLR_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/JKF2D",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_J_CLK_negedge or Tviol_K_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => DFM3_Q_tab,
        DataIn => (
               CLK_ipd, K_delayed, J_delayed, Q_zd, CLK_delayed, CLR_ipd));
      Q_zd := Violation XOR Q_zd;
      J_delayed := J_ipd;
      K_delayed := K_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_JKF2D_VITAL of JKF2D is
   for VITAL_ACT
   end for;
end CFG_JKF2D_VITAL;


----- CELL MAJ3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MAJ3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MAJ3 : entity is TRUE;
end MAJ3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of MAJ3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((C_ipd) AND (B_ipd)) OR ((B_ipd) AND (A_ipd)) OR ((C_ipd) AND
         (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MAJ3_VITAL of MAJ3 is
   for VITAL_ACT
   end for;
end CFG_MAJ3_VITAL;


----- CELL MX2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MX2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MX2 : entity is TRUE;
end MX2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of MX2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := VitalMUX
                 (data => (B_ipd, A_ipd),
                  dselect => (0 => S_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MX2_VITAL of MX2 is
   for VITAL_ACT
   end for;
end CFG_MX2_VITAL;


----- CELL MX2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MX2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MX2A : entity is TRUE;
end MX2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of MX2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((S_ipd) AND (B_ipd)) OR (((NOT S_ipd)) AND ((NOT A_ipd))) OR ((B_ipd) AND ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MX2A_VITAL of MX2A is
   for VITAL_ACT
   end for;
end CFG_MX2A_VITAL;


----- CELL MX2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MX2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MX2B : entity is TRUE;
end MX2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of MX2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((S_ipd) AND ((NOT B_ipd))) OR (((NOT S_ipd)) AND (A_ipd)) OR ((A_ipd) AND ((NOT B_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MX2B_VITAL of MX2B is
   for VITAL_ACT
   end for;
end CFG_MX2B_VITAL;


----- CELL MX2C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MX2C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MX2C : entity is TRUE;
end MX2C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of MX2C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := VitalMUX
                 (data => (B_ipd, A_ipd),
                  dselect => (0 => S_ipd));
      Y_zd := NOT Y_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MX2C_VITAL of MX2C is
   for VITAL_ACT
   end for;
end CFG_MX2C_VITAL;


----- CELL MX4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MX4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0                             :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MX4 : entity is TRUE;
end MX4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of MX4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0_ipd, S0, tipd_S0);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := VitalMUX
                 (data => (D3_ipd, D2_ipd, D1_ipd, D0_ipd),
                  dselect => (S1_ipd, S0_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S1_ipd'last_event, tpd_S1_Y, TRUE),
                 1 => (S0_ipd'last_event, tpd_S0_Y, TRUE),
                 2 => (D3_ipd'last_event, tpd_D3_Y, TRUE),
                 3 => (D2_ipd'last_event, tpd_D2_Y, TRUE),
                 4 => (D1_ipd'last_event, tpd_D1_Y, TRUE),
                 5 => (D0_ipd'last_event, tpd_D0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MX4_VITAL of MX4 is
   for VITAL_ACT
   end for;
end CFG_MX4_VITAL;


----- CELL MXC1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MXC1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      S                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MXC1 : entity is TRUE;
end MXC1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of MXC1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (S_ipd, S, tipd_S);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, S_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   VARIABLE MUX_Out : std_ulogic;

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      --Y_zd :=
      -- ((D_ipd) AND (((B_ipd) AND (S_ipd)) OR ((A_ipd) AND ((NOT S_ipd)))))
      --   OR ((C_ipd) AND ((NOT (((B_ipd) AND (S_ipd)) OR ((A_ipd) AND ((NOT
      --   S_ipd)))))));
      MUX_Out := VitalMUX2(B_ipd, A_ipd, S_ipd);
      Y_zd := VitalMUX2(D_ipd, C_ipd, MUX_Out);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S_ipd'last_event, tpd_S_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MXC1_VITAL of MXC1 is
   for VITAL_ACT
   end for;
end CFG_MXC1_VITAL;


----- CELL MXT -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity MXT is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_S1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0B_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_S0A_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D3_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D2_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D1_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D0_Y                       :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D0                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D2                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D3                        :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0A                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S0B                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_S1                        :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D0                             :	in    STD_ULOGIC;
      D1                             :	in    STD_ULOGIC;
      D2                             :	in    STD_ULOGIC;
      D3                             :	in    STD_ULOGIC;
      S0A                            :	in    STD_ULOGIC;
      S0B                            :	in    STD_ULOGIC;
      S1                             :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of MXT : entity is TRUE;
end MXT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of MXT is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D0_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D1_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D2_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D3_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S0B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL S1_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D0_ipd, D0, tipd_D0);
   VitalWireDelay (D1_ipd, D1, tipd_D1);
   VitalWireDelay (D2_ipd, D2, tipd_D2);
   VitalWireDelay (D3_ipd, D3, tipd_D3);
   VitalWireDelay (S0A_ipd, S0A, tipd_S0A);
   VitalWireDelay (S0B_ipd, S0B, tipd_S0B);
   VitalWireDelay (S1_ipd, S1, tipd_S1);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D0_ipd, D1_ipd, D2_ipd, D3_ipd, S0A_ipd, S0B_ipd, S1_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);
   VARIABLE MUX1_Out, MUX2_Out : std_ulogic;

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      --Y_zd :=
      -- ((S0A_ipd) AND ((NOT S1_ipd)) AND (D1_ipd)) OR (((NOT S0A_ipd)) AND
      --   ((NOT S1_ipd)) AND (D0_ipd)) OR (((NOT S0B_ipd)) AND (S1_ipd) AND
      --   (D2_ipd)) OR ((S0B_ipd) AND (S1_ipd) AND (D3_ipd));
      MUX1_Out := VitalMUX2(D1_ipd, D0_ipd, S0A_ipd);
      MUX2_Out := VitalMUX2(D3_ipd, D2_ipd, S0B_ipd);
      Y_zd := VitalMUX2(MUX2_Out, MUX1_Out, S1_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (S1_ipd'last_event, tpd_S1_Y, TRUE),
                 1 => (S0B_ipd'last_event, tpd_S0B_Y, TRUE),
                 2 => (S0A_ipd'last_event, tpd_S0A_Y, TRUE),
                 3 => (D3_ipd'last_event, tpd_D3_Y, TRUE),
                 4 => (D2_ipd'last_event, tpd_D2_Y, TRUE),
                 5 => (D1_ipd'last_event, tpd_D1_Y, TRUE),
                 6 => (D0_ipd'last_event, tpd_D0_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_MXT_VITAL of MXT is
   for VITAL_ACT
   end for;
end CFG_MXT_VITAL;


----- CELL NAND2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND2 : entity is TRUE;
end NAND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NAND2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) AND (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND2_VITAL of NAND2 is
   for VITAL_ACT
   end for;
end CFG_NAND2_VITAL;


----- CELL NAND2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND2A : entity is TRUE;
end NAND2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NAND2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) AND ((NOT A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND2A_VITAL of NAND2A is
   for VITAL_ACT
   end for;
end CFG_NAND2A_VITAL;


----- CELL NAND2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND2B : entity is TRUE;
end NAND2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NAND2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT B_ipd)) AND ((NOT A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND2B_VITAL of NAND2B is
   for VITAL_ACT
   end for;
end CFG_NAND2B_VITAL;


----- CELL NAND3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND3 : entity is TRUE;
end NAND3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NAND3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) AND (A_ipd) AND (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND3_VITAL of NAND3 is
   for VITAL_ACT
   end for;
end CFG_NAND3_VITAL;


----- CELL NAND3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND3A : entity is TRUE;
end NAND3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NAND3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) AND ((NOT A_ipd)) AND (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND3A_VITAL of NAND3A is
   for VITAL_ACT
   end for;
end CFG_NAND3A_VITAL;


----- CELL NAND3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND3B : entity is TRUE;
end NAND3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NAND3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT B_ipd)) AND ((NOT A_ipd)) AND (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND3B_VITAL of NAND3B is
   for VITAL_ACT
   end for;
end CFG_NAND3B_VITAL;


----- CELL NAND3C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND3C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND3C : entity is TRUE;
end NAND3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NAND3C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND3C_VITAL of NAND3C is
   for VITAL_ACT
   end for;
end CFG_NAND3C_VITAL;


----- CELL NAND4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND4 : entity is TRUE;
end NAND4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NAND4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) AND (A_ipd) AND (C_ipd) AND (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND4_VITAL of NAND4 is
   for VITAL_ACT
   end for;
end CFG_NAND4_VITAL;


----- CELL NAND4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND4A : entity is TRUE;
end NAND4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NAND4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) AND ((NOT A_ipd)) AND (C_ipd) AND (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND4A_VITAL of NAND4A is
   for VITAL_ACT
   end for;
end CFG_NAND4A_VITAL;


----- CELL NAND4B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND4B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND4B : entity is TRUE;
end NAND4B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NAND4B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) AND ((NOT A_ipd)) AND (C_ipd) AND (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND4B_VITAL of NAND4B is
   for VITAL_ACT
   end for;
end CFG_NAND4B_VITAL;


----- CELL NAND4C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND4C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND4C : entity is TRUE;
end NAND4C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NAND4C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd)) AND (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND4C_VITAL of NAND4C is
   for VITAL_ACT
   end for;
end CFG_NAND4C_VITAL;


----- CELL NAND4D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND4D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND4D : entity is TRUE;
end NAND4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NAND4D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd)) AND ((NOT
         D_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND4D_VITAL of NAND4D is
   for VITAL_ACT
   end for;
end CFG_NAND4D_VITAL;


----- CELL NAND5C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NAND5C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NAND5C : entity is TRUE;
end NAND5C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NAND5C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) AND ((NOT A_ipd)) AND ((NOT C_ipd)) AND (D_ipd)
         AND (E_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 4 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NAND5C_VITAL of NAND5C is
   for VITAL_ACT
   end for;
end CFG_NAND5C_VITAL;


----- CELL NOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR2 : entity is TRUE;
end NOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NOR2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) OR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR2_VITAL of NOR2 is
   for VITAL_ACT
   end for;
end CFG_NOR2_VITAL;


----- CELL NOR2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR2A : entity is TRUE;
end NOR2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NOR2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) OR ((NOT A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR2A_VITAL of NOR2A is
   for VITAL_ACT
   end for;
end CFG_NOR2A_VITAL;


----- CELL NOR2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR2B : entity is TRUE;
end NOR2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NOR2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT B_ipd)) OR ((NOT A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR2B_VITAL of NOR2B is
   for VITAL_ACT
   end for;
end CFG_NOR2B_VITAL;


----- CELL NOR3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR3 : entity is TRUE;
end NOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NOR3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) OR (A_ipd) OR (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR3_VITAL of NOR3 is
   for VITAL_ACT
   end for;
end CFG_NOR3_VITAL;


----- CELL NOR3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR3A : entity is TRUE;
end NOR3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NOR3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) OR ((NOT A_ipd)) OR (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR3A_VITAL of NOR3A is
   for VITAL_ACT
   end for;
end CFG_NOR3A_VITAL;


----- CELL NOR3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR3B : entity is TRUE;
end NOR3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NOR3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT B_ipd)) OR ((NOT A_ipd)) OR (C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR3B_VITAL of NOR3B is
   for VITAL_ACT
   end for;
end CFG_NOR3B_VITAL;


----- CELL NOR3C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR3C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR3C : entity is TRUE;
end NOR3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NOR3C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT B_ipd)) OR ((NOT A_ipd)) OR ((NOT C_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR3C_VITAL of NOR3C is
   for VITAL_ACT
   end for;
end CFG_NOR3C_VITAL;


----- CELL NOR4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR4 : entity is TRUE;
end NOR4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NOR4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) OR (A_ipd) OR (C_ipd) OR (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR4_VITAL of NOR4 is
   for VITAL_ACT
   end for;
end CFG_NOR4_VITAL;


----- CELL NOR4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR4A : entity is TRUE;
end NOR4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NOR4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) OR ((NOT A_ipd)) OR (C_ipd) OR (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR4A_VITAL of NOR4A is
   for VITAL_ACT
   end for;
end CFG_NOR4A_VITAL;


----- CELL NOR4B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR4B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR4B : entity is TRUE;
end NOR4B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NOR4B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) OR ((NOT A_ipd)) OR (C_ipd) OR (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR4B_VITAL of NOR4B is
   for VITAL_ACT
   end for;
end CFG_NOR4B_VITAL;


----- CELL NOR4C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR4C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR4C : entity is TRUE;
end NOR4C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NOR4C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) OR ((NOT A_ipd)) OR ((NOT C_ipd)) OR (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR4C_VITAL of NOR4C is
   for VITAL_ACT
   end for;
end CFG_NOR4C_VITAL;


----- CELL NOR4D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR4D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR4D : entity is TRUE;
end NOR4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NOR4D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) OR ((NOT A_ipd)) OR ((NOT C_ipd)) OR ((NOT
         D_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR4D_VITAL of NOR4D is
   for VITAL_ACT
   end for;
end CFG_NOR4D_VITAL;


----- CELL NOR5C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity NOR5C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of NOR5C : entity is TRUE;
end NOR5C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of NOR5C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT B_ipd)) OR ((NOT A_ipd)) OR ((NOT C_ipd)) OR (D_ipd) OR
         (E_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 4 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_NOR5C_VITAL of NOR5C is
   for VITAL_ACT
   end for;
end CFG_NOR5C_VITAL;


----- CELL OA1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA1 : entity is TRUE;
end OA1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OA1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) AND ((B_ipd) OR (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA1_VITAL of OA1 is
   for VITAL_ACT
   end for;
end CFG_OA1_VITAL;


----- CELL OA1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA1A : entity is TRUE;
end OA1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OA1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) AND ((B_ipd) OR ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA1A_VITAL of OA1A is
   for VITAL_ACT
   end for;
end CFG_OA1A_VITAL;


----- CELL OA1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA1B : entity is TRUE;
end OA1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OA1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) AND ((B_ipd) OR (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA1B_VITAL of OA1B is
   for VITAL_ACT
   end for;
end CFG_OA1B_VITAL;


----- CELL OA1C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA1C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA1C : entity is TRUE;
end OA1C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OA1C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) AND ((B_ipd) OR ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA1C_VITAL of OA1C is
   for VITAL_ACT
   end for;
end CFG_OA1C_VITAL;


----- CELL OA2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA2 : entity is TRUE;
end OA2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OA2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((D_ipd) OR (C_ipd)) AND ((B_ipd) OR (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA2_VITAL of OA2 is
   for VITAL_ACT
   end for;
end CFG_OA2_VITAL;


----- CELL OA2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA2A : entity is TRUE;
end OA2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OA2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((D_ipd) OR (C_ipd)) AND ((B_ipd) OR ((NOT A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA2A_VITAL of OA2A is
   for VITAL_ACT
   end for;
end CFG_OA2A_VITAL;


----- CELL OA3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA3 : entity is TRUE;
end OA3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OA3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) AND ((B_ipd) OR (A_ipd)) AND (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA3_VITAL of OA3 is
   for VITAL_ACT
   end for;
end CFG_OA3_VITAL;


----- CELL OA3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA3A : entity is TRUE;
end OA3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OA3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) AND ((B_ipd) OR (A_ipd)) AND (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA3A_VITAL of OA3A is
   for VITAL_ACT
   end for;
end CFG_OA3A_VITAL;


----- CELL OA3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA3B : entity is TRUE;
end OA3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OA3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT C_ipd)) AND ((B_ipd) OR ((NOT A_ipd))) AND (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA3B_VITAL of OA3B is
   for VITAL_ACT
   end for;
end CFG_OA3B_VITAL;


----- CELL OA4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA4 : entity is TRUE;
end OA4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OA4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (D_ipd) AND ((B_ipd) OR (A_ipd) OR (C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA4_VITAL of OA4 is
   for VITAL_ACT
   end for;
end CFG_OA4_VITAL;


----- CELL OA4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA4A : entity is TRUE;
end OA4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OA4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (D_ipd) AND ((B_ipd) OR (A_ipd) OR ((NOT C_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA4A_VITAL of OA4A is
   for VITAL_ACT
   end for;
end CFG_OA4A_VITAL;


----- CELL OA5 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OA5 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OA5 : entity is TRUE;
end OA5;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OA5 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((D_ipd) OR (A_ipd)) AND ((B_ipd) OR (A_ipd) OR (C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OA5_VITAL of OA5 is
   for VITAL_ACT
   end for;
end CFG_OA5_VITAL;


----- CELL OAI1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI1 : entity is TRUE;
end OAI1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OAI1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((C_ipd) AND ((B_ipd) OR (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OAI1_VITAL of OAI1 is
   for VITAL_ACT
   end for;
end CFG_OAI1_VITAL;


----- CELL OAI2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI2A : entity is TRUE;
end OAI2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OAI2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT (((NOT D_ipd)) AND ((B_ipd) OR (A_ipd) OR (C_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OAI2A_VITAL of OAI2A is
   for VITAL_ACT
   end for;
end CFG_OAI2A_VITAL;


----- CELL OAI3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI3 : entity is TRUE;
end OAI3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OAI3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((C_ipd) AND ((B_ipd) OR (A_ipd)) AND (D_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OAI3_VITAL of OAI3 is
   for VITAL_ACT
   end for;
end CFG_OAI3_VITAL;


----- CELL OAI3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OAI3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OAI3A : entity is TRUE;
end OAI3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OAI3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       (NOT (((NOT C_ipd)) AND ((B_ipd) OR (A_ipd)) AND ((NOT D_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 3 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OAI3A_VITAL of OAI3A is
   for VITAL_ACT
   end for;
end CFG_OAI3A_VITAL;


----- CELL OBDLHS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OBDLHS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OBDLHS : entity is TRUE;
end OBDLHS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OBDLHS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_PAD : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/OBDLHS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/OBDLHS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Pviol_G;
      VitalStateTable(
        Result => PAD_zd,
        PreviousDataIn => PrevData_PAD,
        StateTable => DL1_Q_tab,
        DataIn => (
               D_ipd, G_ipd));
      PAD_zd := Violation XOR PAD_zd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_PAD, TRUE),
                 1 => (G_ipd'last_event, tpd_G_PAD, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OBDLHS_VITAL of OBDLHS is
   for VITAL_ACT
   end for;
end CFG_OBDLHS_VITAL;


----- CELL OBHS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OBHS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OBHS : entity is TRUE;
end OBHS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OBHS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := TO_X01(D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_PAD, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OBHS_VITAL of OBHS is
   for VITAL_ACT
   end for;
end CFG_OBHS_VITAL;


----- CELL OR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR2 : entity is TRUE;
end OR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OR2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) OR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR2_VITAL of OR2 is
   for VITAL_ACT
   end for;
end CFG_OR2_VITAL;


----- CELL OR2A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR2A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR2A : entity is TRUE;
end OR2A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OR2A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) OR ((NOT A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR2A_VITAL of OR2A is
   for VITAL_ACT
   end for;
end CFG_OR2A_VITAL;


----- CELL OR2B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR2B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR2B : entity is TRUE;
end OR2B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OR2B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) OR ((NOT A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR2B_VITAL of OR2B is
   for VITAL_ACT
   end for;
end CFG_OR2B_VITAL;


----- CELL OR3 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR3 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR3 : entity is TRUE;
end OR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OR3 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) OR (A_ipd) OR (C_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR3_VITAL of OR3 is
   for VITAL_ACT
   end for;
end CFG_OR3_VITAL;


----- CELL OR3A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR3A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR3A : entity is TRUE;
end OR3A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OR3A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) OR ((NOT A_ipd)) OR (C_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR3A_VITAL of OR3A is
   for VITAL_ACT
   end for;
end CFG_OR3A_VITAL;


----- CELL OR3B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR3B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR3B : entity is TRUE;
end OR3B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OR3B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) OR ((NOT A_ipd)) OR (C_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR3B_VITAL of OR3B is
   for VITAL_ACT
   end for;
end CFG_OR3B_VITAL;


----- CELL OR3C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR3C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR3C : entity is TRUE;
end OR3C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OR3C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) OR ((NOT A_ipd)) OR ((NOT C_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR3C_VITAL of OR3C is
   for VITAL_ACT
   end for;
end CFG_OR3C_VITAL;


----- CELL OR4 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR4 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR4 : entity is TRUE;
end OR4;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OR4 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) OR (A_ipd) OR (C_ipd) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR4_VITAL of OR4 is
   for VITAL_ACT
   end for;
end CFG_OR4_VITAL;


----- CELL OR4A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR4A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR4A : entity is TRUE;
end OR4A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OR4A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) OR ((NOT A_ipd)) OR (C_ipd) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 1 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 3 => (B_ipd'last_event, tpd_B_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR4A_VITAL of OR4A is
   for VITAL_ACT
   end for;
end CFG_OR4A_VITAL;


----- CELL OR4B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR4B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR4B : entity is TRUE;
end OR4B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OR4B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) OR ((NOT A_ipd)) OR (C_ipd) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 3 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR4B_VITAL of OR4B is
   for VITAL_ACT
   end for;
end CFG_OR4B_VITAL;


----- CELL OR4C -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR4C is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR4C : entity is TRUE;
end OR4C;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OR4C is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := ((NOT B_ipd)) OR ((NOT A_ipd)) OR ((NOT C_ipd)) OR (D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 1 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 2 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR4C_VITAL of OR4C is
   for VITAL_ACT
   end for;
end CFG_OR4C_VITAL;


----- CELL OR4D -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR4D is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR4D : entity is TRUE;
end OR4D;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OR4D is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((NOT B_ipd)) OR ((NOT A_ipd)) OR ((NOT C_ipd)) OR ((NOT D_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 1 => (C_ipd'last_event, tpd_C_Y, TRUE),
                 2 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 3 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR4D_VITAL of OR4D is
   for VITAL_ACT
   end for;
end CFG_OR4D_VITAL;


----- CELL OR5B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OR5B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_D_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OR5B : entity is TRUE;
end OR5B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OR5B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';
   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd, D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd :=
       ((NOT B_ipd)) OR ((NOT A_ipd)) OR (C_ipd) OR (D_ipd) OR (E_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (E_ipd'last_event, tpd_E_Y, TRUE),
                 3 => (D_ipd'last_event, tpd_D_Y, TRUE),
                 4 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OR5B_VITAL of OR5B is
   for VITAL_ACT
   end for;
end CFG_OR5B_VITAL;


----- CELL ORH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity ORH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of ORH : entity is TRUE;
end ORH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of ORH is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_PAD : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/ORH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/ORH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => PAD_zd,
        PreviousDataIn => PrevData_PAD,
        StateTable => DF1_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd));
      PAD_zd := Violation XOR PAD_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_PAD, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_ORH_VITAL of ORH is
   for VITAL_ACT
   end for;
end CFG_ORH_VITAL;


----- CELL ORIH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity ORIH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of ORIH : entity is TRUE;
end ORIH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of ORIH is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_PAD : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/ORIH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/ORIH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => PAD_zd,
        PreviousDataIn => PrevData_PAD,
        StateTable => DF1A_QN_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd));
      PAD_zd := Violation XOR PAD_zd;
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (CLK_ipd'last_event, tpd_CLK_PAD, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_ORIH_VITAL of ORIH is
   for VITAL_ACT
   end for;
end CFG_ORIH_VITAL;


----- CELL ORITH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity ORITH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of ORITH : entity is TRUE;
end ORITH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of ORITH is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_PAD : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zdi : STD_LOGIC is Results(1);
   VARIABLE PAD_zd : STD_ULOGIC := 'X';

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/ORITH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/ORITH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => PAD_zdi,
        PreviousDataIn => PrevData_PAD,
        StateTable => DF1A_QN_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd));
      PAD_zdi := Violation XOR PAD_zdi;
      PAD_zd := VitalBUFIF0 (data => PAD_zdi,
             enable => (NOT E_ipd));
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_PAD, TRUE),
                 1 => (CLK_ipd'last_event, VitalExtendToFillDelay(tpd_CLK_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_ORITH_VITAL of ORITH is
   for VITAL_ACT
   end for;
end CFG_ORITH_VITAL;


----- CELL ORTH -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity ORTH is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_CLK_PAD                    :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_D_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_D_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of ORTH : entity is TRUE;
end ORTH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of ORTH is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, CLK_ipd)

   -- timing check results
   VARIABLE Tviol_D_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_PAD : STD_LOGIC_VECTOR(0 to 2);
   VARIABLE D_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zdi : STD_LOGIC is Results(1);
   VARIABLE PAD_zd : STD_ULOGIC := 'X';

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_CLK_posedge,
          TimingData              => Tmkr_D_CLK_posedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_CLK_noedge_posedge,
          SetupLow                => tsetup_D_CLK_noedge_posedge,
          HoldHigh                => thold_D_CLK_noedge_posedge,
          HoldLow                 => thold_D_CLK_noedge_posedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/ORTH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/ORTH",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_CLK_posedge or Pviol_CLK;
      VitalStateTable(
        Result => PAD_zdi,
        PreviousDataIn => PrevData_PAD,
        StateTable => DF1_Q_tab,
        DataIn => (
               CLK_delayed, D_delayed, CLK_ipd));
      PAD_zdi := Violation XOR PAD_zdi;
      PAD_zd := VitalBUFIF0 (data => PAD_zdi,
             enable => (NOT E_ipd));
      D_delayed := D_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_PAD, TRUE),
                 1 => (CLK_ipd'last_event, VitalExtendToFillDelay(tpd_CLK_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_ORTH_VITAL of ORTH is
   for VITAL_ACT
   end for;
end CFG_ORTH_VITAL;


----- CELL OUTBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity OUTBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of OUTBUF : entity is TRUE;
end OUTBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of OUTBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := TO_X01(D_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (D_ipd'last_event, tpd_D_PAD, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_OUTBUF_VITAL of OUTBUF is
   for VITAL_ACT
   end for;
end CFG_OUTBUF_VITAL;


----- CELL QCLKBUF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity QCLKBUF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_PAD_Y                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_PAD                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      PAD                            :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of QCLKBUF : entity is TRUE;
end QCLKBUF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of QCLKBUF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL PAD_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (PAD_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(PAD_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (PAD_ipd'last_event, tpd_PAD_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_QCLKBUF_VITAL of QCLKBUF is
   for VITAL_ACT
   end for;
end CFG_QCLKBUF_VITAL;


----- CELL QCLKINT -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity QCLKINT is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of QCLKINT : entity is TRUE;
end QCLKINT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of QCLKINT is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := TO_X01(A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_QCLKINT_VITAL of QCLKINT is
   for VITAL_ACT
   end for;
end CFG_QCLKINT_VITAL;


























-----------------------------------------------------------------
--  Proxy Modeling, Inc. 
--
--  Actel RAM4FA VHDL behavioral model
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - Jan/22/96 - Initial Delivery
-- 1.1 - 12/6/96 by DNW - Modified SL_TO_INT.
-- 1.2 - 3/3/97 by DNW - WDx_delayed variables added.
-- 1.3 - 3/6/98 by DNW - Issue "unknown" msg. only if 0/1->X Xtion.
-- 1.4 - 5/27/98 by DNW - Initaialize _ipd signals to X instead of 0.
-- 
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity RAM4FA is
  GENERIC (
        tipd_RDAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RDAD5_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD5_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD5_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD5_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_WRAD5_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of RAM4FA : entity is TRUE;
  
end RAM4FA;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM4FA is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal WRAD5_ipd : std_ulogic := 'X';
  signal WRAD4_ipd : std_ulogic := 'X';
  signal WRAD3_ipd : std_ulogic := 'X';
  signal WRAD2_ipd : std_ulogic := 'X';
  signal WRAD1_ipd : std_ulogic := 'X';
  signal WRAD0_ipd : std_ulogic := 'X';
  signal WD3_ipd : std_ulogic := 'X';
  signal WD2_ipd : std_ulogic := 'X';
  signal WD1_ipd : std_ulogic := 'X';
  signal WD0_ipd : std_ulogic := 'X';
  signal RDAD5_ipd : std_ulogic := 'X';
  signal RDAD4_ipd : std_ulogic := 'X';
  signal RDAD3_ipd : std_ulogic := 'X';
  signal RDAD2_ipd : std_ulogic := 'X';
  signal RDAD1_ipd : std_ulogic := 'X';
  signal RDAD0_ipd : std_ulogic := 'X';
  signal BLKEN_ipd : std_ulogic := 'X';
  signal WEN_ipd : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  type MEM is array(0 to 63) of std_ulogic_vector(3 downto 0);
   signal RAM_TMP : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (WRAD5_ipd, WRAD5, VitalExtendToFillDelay(tipd_WRAD5));
    VitalWireDelay (WRAD4_ipd, WRAD4, VitalExtendToFillDelay(tipd_WRAD4));
    VitalWireDelay (WRAD3_ipd, WRAD3, VitalExtendToFillDelay(tipd_WRAD3));
    VitalWireDelay (WRAD2_ipd, WRAD2, VitalExtendToFillDelay(tipd_WRAD2));
    VitalWireDelay (WRAD1_ipd, WRAD1, VitalExtendToFillDelay(tipd_WRAD1));
    VitalWireDelay (WRAD0_ipd, WRAD0, VitalExtendToFillDelay(tipd_WRAD0));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (RDAD5_ipd, RDAD5, VitalExtendToFillDelay(tipd_RDAD5));
    VitalWireDelay (RDAD4_ipd, RDAD4, VitalExtendToFillDelay(tipd_RDAD4));
    VitalWireDelay (RDAD3_ipd, RDAD3, VitalExtendToFillDelay(tipd_RDAD3));
    VitalWireDelay (RDAD2_ipd, RDAD2, VitalExtendToFillDelay(tipd_RDAD2));
    VitalWireDelay (RDAD1_ipd, RDAD1, VitalExtendToFillDelay(tipd_RDAD1));
    VitalWireDelay (RDAD0_ipd, RDAD0, VitalExtendToFillDelay(tipd_RDAD0));
    VitalWireDelay (BLKEN_ipd, BLKEN, VitalExtendToFillDelay(tipd_BLKEN));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (RDAD5_ipd, RDAD4_ipd, RDAD3_ipd, RDAD2_ipd, 
		RDAD1_ipd, RDAD0_ipd, 
		WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd, WRAD5_ipd, WRAD4_ipd, 
		WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, WEN_ipd, 
		BLKEN_ipd, BLKENS, WCLK_ipd, RAM_TMP)

     --  Write Timing Check Results
     variable Tviol_WD3_WCLK_negedge : X01 := '0';
     variable TmDt_WD3_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_negedge : X01 := '0';
     variable TmDt_WD2_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_negedge : X01 := '0';
     variable TmDt_WD1_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_negedge : X01 := '0';
     variable TmDt_WD0_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD5_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD5_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD4_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD4_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD3_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD3_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD2_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD2_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD1_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD1_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD0_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD0_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_negedge : X01 := '0';
     variable TmDt_WEN_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_BLKEN_WCLK_negedge : X01 := '0';
     variable TmDt_BLKEN_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     --type SL_TO_INT is array(std_ulogic range <>) of integer;
     --constant INT :SL_TO_INT('U' to '-') := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;
  
     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable WEN_delayed : std_ulogic := 'X';
     variable WEN_previous : std_ulogic := 'X';
     variable BLKEN_delayed : std_ulogic := 'X';
     variable BLKEN_previous : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WRAD5_delayed : std_ulogic := 'X';
     variable WRAD4_delayed : std_ulogic := 'X';
     variable WRAD3_delayed : std_ulogic := 'X';
     variable WRAD2_delayed : std_ulogic := 'X';
     variable WRAD1_delayed : std_ulogic := 'X';
     variable WRAD0_delayed : std_ulogic := 'X';
     variable WRAD5_previous : std_ulogic := 'X';
     variable WRAD4_previous : std_ulogic := 'X';
     variable WRAD3_previous : std_ulogic := 'X';
     variable WRAD2_previous : std_ulogic := 'X';
     variable WRAD1_previous : std_ulogic := 'X';
     variable WRAD0_previous : std_ulogic := 'X';
     variable RDAD5_previous : std_ulogic := 'X';
     variable RDAD4_previous : std_ulogic := 'X';
     variable RDAD3_previous : std_ulogic := 'X';
     variable RDAD2_previous : std_ulogic := 'X';
     variable RDAD1_previous : std_ulogic := 'X';
     variable RDAD0_previous : std_ulogic := 'X';
  
  begin  --  process VITALBehavior 

    if (TimingCheckOn) then

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup BLKEN high or low before WCLK falling
      --   Hold  BLKEN high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_BLKEN_WCLK_negedge,
                            TmDt_BLKEN_WCLK_negedge,
                            BLKEN_ipd, "BLKEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_BLKEN_WCLK_noedge_negedge,
                            tsetup_BLKEN_WCLK_noedge_negedge,
                            thold_BLKEN_WCLK_noedge_negedge,
                            thold_BLKEN_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WRAD high or low before WCLK falling
      --   Hold  WRAD high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_WRAD5_WCLK_negedge,
                            TmDt_WRAD5_WCLK_negedge,
                            WRAD5_ipd, "WRAD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD5_WCLK_noedge_negedge,
                            tsetup_WRAD5_WCLK_noedge_negedge,
                            thold_WRAD5_WCLK_noedge_negedge,
                            thold_WRAD5_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD4_WCLK_negedge,
                            TmDt_WRAD4_WCLK_negedge,
                            WRAD4_ipd, "WRAD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD4_WCLK_noedge_negedge,
                            tsetup_WRAD4_WCLK_noedge_negedge,
                            thold_WRAD4_WCLK_noedge_negedge,
                            thold_WRAD4_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD3_WCLK_negedge,
                            TmDt_WRAD3_WCLK_negedge,
                            WRAD3_ipd, "WRAD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD3_WCLK_noedge_negedge,
                            tsetup_WRAD3_WCLK_noedge_negedge,
                            thold_WRAD3_WCLK_noedge_negedge,
                            thold_WRAD3_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD2_WCLK_negedge,
                            TmDt_WRAD2_WCLK_negedge,
                            WRAD2_ipd, "WRAD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD2_WCLK_noedge_negedge,
                            tsetup_WRAD2_WCLK_noedge_negedge,
                            thold_WRAD2_WCLK_noedge_negedge,
                            thold_WRAD2_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD1_WCLK_negedge,
                            TmDt_WRAD1_WCLK_negedge,
                            WRAD1_ipd, "WRAD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD1_WCLK_noedge_negedge,
                            tsetup_WRAD1_WCLK_noedge_negedge,
                            thold_WRAD1_WCLK_noedge_negedge,
                            thold_WRAD1_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD0_WCLK_negedge,
                            TmDt_WRAD0_WCLK_negedge,
                            WRAD0_ipd, "WRAD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD0_WCLK_noedge_negedge,
                            tsetup_WRAD0_WCLK_noedge_negedge,
                            thold_WRAD0_WCLK_noedge_negedge,
                            thold_WRAD0_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WD high or low before WCLK falling
      --   Hold  WD high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_negedge,
                            TmDt_WD3_WCLK_negedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_noedge_negedge,
                            tsetup_WD3_WCLK_noedge_negedge,
                            thold_WD3_WCLK_noedge_negedge,
                            thold_WD3_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_negedge,
                            TmDt_WD2_WCLK_negedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_noedge_negedge,
                            tsetup_WD2_WCLK_noedge_negedge,
                            thold_WD2_WCLK_noedge_negedge,
                            thold_WD2_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_negedge,
                            TmDt_WD1_WCLK_negedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_noedge_negedge,
                            tsetup_WD1_WCLK_noedge_negedge,
                            thold_WD1_WCLK_noedge_negedge,
                            thold_WD1_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_negedge,
                            TmDt_WD0_WCLK_negedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_noedge_negedge,
                            tsetup_WD0_WCLK_noedge_negedge,
                            thold_WD0_WCLK_noedge_negedge,
                            thold_WD0_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup WEN high before WCLK falling
      --   Hold  WEN high after WCLK falling

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_negedge,
                            TmDt_WEN_WCLK_negedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_noedge_negedge,
                            tsetup_WEN_WCLK_noedge_negedge,
                            thold_WEN_WCLK_noedge_negedge,
                            thold_WEN_WCLK_noedge_negedge,
                            (To_X01(BLKEN_ipd)=BLKENS),
                            '\',
                            InstancePath & "/RAM4FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM4FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
    
    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      -- Convert Write Address Signal to Integer
      WADDR := ((INT(WRAD5_delayed)*32)+(INT(WRAD4_delayed)*16)+(INT(WRAD3_delayed)*8)+
		(INT(WRAD2_delayed)*4)+(INT(WRAD1_delayed)*2)+(INT(WRAD0_delayed)));

      if (TO_X01(WCLK_ipd)='X') then
        if (TO_X01(WCLK_previous) /= 'X') then
	  assert false
	  report ": WCLK unknown"
	  severity Warning;
	end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='0')) then
	case TO_X01(WEN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (TO_X01(BLKEN_delayed) = 'X') then
              if (TO_X01(BLKEN_previous) /= 'X') then
	        assert false
	        report ": BLKEN unknown"
	        severity Warning;
	      end if;
	    elsif (TO_X01(BLKEN_delayed) = BLKENS) then
	      if (WADDR < 0) then
		if (TO_X01(WRAD5_delayed) = 'X') and (TO_X01(WRAD5_previous) /= 'X') then
		  assert false
		  report ": WRAD5 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD4_delayed) = 'X') and (TO_X01(WRAD4_previous) /= 'X') then
		  assert false
		  report ": WRAD4 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD3_delayed) = 'X') and (TO_X01(WRAD3_previous) /= 'X') then
		  assert false
		  report ": WRAD3 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD2_delayed) = 'X') and (TO_X01(WRAD2_previous) /= 'X') then
		  assert false
		  report ": WRAD2 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD1_delayed) = 'X') and (TO_X01(WRAD1_previous) /= 'X') then
		  assert false
		  report ": WRAD1 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD0_delayed) = 'X') and (TO_X01(WRAD0_previous) /= 'X') then
		  assert false
		  report ": WRAD0 unknown"
		  severity Warning;
		end if;
	      else 
		RAM_TMP(WADDR) <= WD3_delayed & WD2_delayed & WD1_delayed & WD0_delayed ; 
	      end if;
	    else
	      null;
	    end if;
	  when others =>
            if (TO_X01(WEN_previous) /= 'X') then
	      assert false
	      report ": WEN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      -- Convert Read Address Signal to Integer
      RADDR := ((INT(RDAD5_ipd)*32)+(INT(RDAD4_ipd)*16)+(INT(RDAD3_ipd)*8)+
		(INT(RDAD2_ipd)*4)+(INT(RDAD1_ipd)*2)+(INT(RDAD0_ipd)));

      if (RADDR < 0) then
	RD3_zd := 'X';
	RD2_zd := 'X';
	RD1_zd := 'X';
	RD0_zd := 'X';
	if (TO_X01(RDAD5_ipd) = 'X') and (TO_X01(RDAD5_previous) /= 'X') then
          assert false
	  report ": RDAD5 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD4_ipd) = 'X') and (TO_X01(RDAD4_previous) /= 'X') then
	  assert false
	  report ": RDAD4 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD3_ipd) = 'X') and (TO_X01(RDAD3_previous) /= 'X') then
	  assert false
	  report ": RDAD3 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD2_ipd) = 'X') and (TO_X01(RDAD2_previous) /= 'X') then
	  assert false
	  report ": RDAD2 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD1_ipd) = 'X') and (TO_X01(RDAD1_previous) /= 'X') then
	  assert false
	  report ": RDAD1 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD0_ipd) = 'X') and (TO_X01(RDAD0_previous) /= 'X') then
	  assert false
	  report ": RDAD0 unknown"
	  severity Warning;
	end if;
      else
	RD3_zd := RAM_TMP(RADDR)(3);
	RD2_zd := RAM_TMP(RADDR)(2);
	RD1_zd := RAM_TMP(RADDR)(1);
	RD0_zd := RAM_TMP(RADDR)(0);
      end if;
      
      WCLK_previous := WCLK_ipd;
      WEN_previous := WEN_delayed;
      WEN_delayed := WEN_ipd;
      BLKEN_previous := BLKEN_delayed;
      BLKEN_delayed := BLKEN_ipd;
      WD3_delayed := WD3_ipd;
      WD2_delayed := WD2_ipd;
      WD1_delayed := WD1_ipd;
      WD0_delayed := WD0_ipd;
      WRAD5_previous := WRAD5_delayed;
      WRAD4_previous := WRAD4_delayed;
      WRAD3_previous := WRAD3_delayed;
      WRAD2_previous := WRAD2_delayed;
      WRAD1_previous := WRAD1_delayed;
      WRAD0_previous := WRAD0_delayed;
      WRAD5_delayed := WRAD5_ipd;
      WRAD4_delayed := WRAD4_ipd;
      WRAD3_delayed := WRAD3_ipd;
      WRAD2_delayed := WRAD2_ipd;
      WRAD1_delayed := WRAD1_ipd;
      WRAD0_delayed := WRAD0_ipd;
      RDAD5_previous := RDAD5_ipd;
      RDAD4_previous := RDAD4_ipd;
      RDAD3_previous := RDAD3_ipd;
      RDAD2_previous := RDAD2_ipd;
      RDAD1_previous := RDAD1_ipd;
      RDAD0_previous := RDAD0_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD3,
	GlitchData => RD3_GlitchData,
	OutSignalName => "RD3",
	OutTemp => RD3_zd,
	Paths => (0 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD3), TRUE),
		  1 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
		  2 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
		  3 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
		  4 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  5 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  6 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD3), TRUE),
                  7 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  8 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  9 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  10 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  11 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  12 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD3), TRUE),
                  13 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  14 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  15 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  16 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  17 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  18 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD3), TRUE),
                  19 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  20 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  21 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  22 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  23 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  24 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD3), TRUE),
                  25 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  26 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  27 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  28 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  29 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  30 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD3), TRUE),
                  31 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  32 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  33 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  34 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  35 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD2,
	GlitchData => RD2_GlitchData,
	OutSignalName => "RD2",
	OutTemp => RD2_zd,
	Paths => (0 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD2), TRUE),
		  1 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
		  2 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
		  3 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
		  4 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  5 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  6 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD2), TRUE),
                  7 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  8 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  9 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  10 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  11 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  12 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD2), TRUE),
                  13 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  14 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  15 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  16 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  17 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  18 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD2), TRUE),
                  19 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  20 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  21 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  22 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  23 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  24 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD2), TRUE),
                  25 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  26 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  27 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  28 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  29 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  30 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD2), TRUE),
                  31 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  32 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  33 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  34 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  35 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD1,
	GlitchData => RD1_GlitchData,
	OutSignalName => "RD1",
	OutTemp => RD1_zd,
	Paths => (0 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD1), TRUE),
		  1 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
		  2 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
		  3 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
		  4 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  5 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  6 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD1), TRUE),
                  7 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  8 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  9 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  10 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  11 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  12 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD1), TRUE),
                  13 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  14 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  15 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  16 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  17 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  18 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD1), TRUE),
                  19 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  20 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  21 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  22 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  23 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  24 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD1), TRUE),
                  25 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  26 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  27 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  28 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  29 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  30 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD1), TRUE),
                  31 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  32 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  33 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  34 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  35 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD0,
	GlitchData => RD0_GlitchData,
	OutSignalName => "RD0",
	OutTemp => RD0_zd,
	Paths => (0 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD0), TRUE),
		  1 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
		  2 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
		  3 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
		  4 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  5 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  6 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD0), TRUE),
                  7 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  8 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  9 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  10 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  11 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  12 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD0), TRUE),
                  13 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  14 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  15 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  16 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  17 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  18 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD0), TRUE),
                  19 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  20 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  21 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  22 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  23 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  24 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD0), TRUE),
                  25 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  26 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  27 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  28 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  29 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  30 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD0), TRUE),
                  31 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  32 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  33 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  34 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  35 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

  end process VITALBehavior;

end VITAL_ACT;
-----------------------------------------------------------------
--  Proxy Modeling, Inc. 
--
--  Actel RAM4FF VHDL behavioral model
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - Jan/22/96 - Initial Delivery
-- 1.1 - 12/6/96 by DNW - Modified SL_TO_INT.
-- 1.2 - 3/3/97 by DNW - WDx_delayed variables added.
-- 1.3 - 3/6/98 by DNW - Issue "unknown" msg. only if 0/1->X Xtion.
-- 1.4 - 5/27/98 by DNW - Initaialize _ipd signals to X instead of 0.
-- 
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity RAM4FF is
  GENERIC (
        tipd_RDAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD5_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of RAM4FF : entity is TRUE;
  
end RAM4FF;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM4FF is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal WRAD5_ipd : std_ulogic := 'X';
  signal WRAD4_ipd : std_ulogic := 'X';
  signal WRAD3_ipd : std_ulogic := 'X';
  signal WRAD2_ipd : std_ulogic := 'X';
  signal WRAD1_ipd : std_ulogic := 'X';
  signal WRAD0_ipd : std_ulogic := 'X';
  signal WD3_ipd : std_ulogic := 'X';
  signal WD2_ipd : std_ulogic := 'X';
  signal WD1_ipd : std_ulogic := 'X';
  signal WD0_ipd : std_ulogic := 'X';
  signal RDAD5_ipd : std_ulogic := 'X';
  signal RDAD4_ipd : std_ulogic := 'X';
  signal RDAD3_ipd : std_ulogic := 'X';
  signal RDAD2_ipd : std_ulogic := 'X';
  signal RDAD1_ipd : std_ulogic := 'X';
  signal RDAD0_ipd : std_ulogic := 'X';
  signal BLKEN_ipd : std_ulogic := 'X';
  signal WEN_ipd : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal REN_ipd : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  type MEM is array(0 to 63) of std_ulogic_vector(3 downto 0);
   signal RAM_TMP : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (WRAD5_ipd, WRAD5, VitalExtendToFillDelay(tipd_WRAD5));
    VitalWireDelay (WRAD4_ipd, WRAD4, VitalExtendToFillDelay(tipd_WRAD4));
    VitalWireDelay (WRAD3_ipd, WRAD3, VitalExtendToFillDelay(tipd_WRAD3));
    VitalWireDelay (WRAD2_ipd, WRAD2, VitalExtendToFillDelay(tipd_WRAD2));
    VitalWireDelay (WRAD1_ipd, WRAD1, VitalExtendToFillDelay(tipd_WRAD1));
    VitalWireDelay (WRAD0_ipd, WRAD0, VitalExtendToFillDelay(tipd_WRAD0));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (RDAD5_ipd, RDAD5, VitalExtendToFillDelay(tipd_RDAD5));
    VitalWireDelay (RDAD4_ipd, RDAD4, VitalExtendToFillDelay(tipd_RDAD4));
    VitalWireDelay (RDAD3_ipd, RDAD3, VitalExtendToFillDelay(tipd_RDAD3));
    VitalWireDelay (RDAD2_ipd, RDAD2, VitalExtendToFillDelay(tipd_RDAD2));
    VitalWireDelay (RDAD1_ipd, RDAD1, VitalExtendToFillDelay(tipd_RDAD1));
    VitalWireDelay (RDAD0_ipd, RDAD0, VitalExtendToFillDelay(tipd_RDAD0));
    VitalWireDelay (BLKEN_ipd, BLKEN, VitalExtendToFillDelay(tipd_BLKEN));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (REN_ipd, REN, VitalExtendToFillDelay(tipd_REN));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (RDAD5_ipd, RDAD4_ipd, RDAD3_ipd, RDAD2_ipd, 
		RDAD1_ipd, RDAD0_ipd, REN_ipd, RCLK_ipd, 
		WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd, WRAD5_ipd, WRAD4_ipd, 
		WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, WEN_ipd, 
		BLKEN_ipd, BLKENS, WCLK_ipd)

     --  Read Timing Check Results
     variable Tviol_RDAD5_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD5_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD4_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD4_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD3_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD3_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD2_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD2_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD1_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD1_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD0_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD0_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_REN_RCLK_negedge : X01 := '0';
     variable TmDt_REN_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_WD3_WCLK_negedge : X01 := '0';
     variable TmDt_WD3_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_negedge : X01 := '0';
     variable TmDt_WD2_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_negedge : X01 := '0';
     variable TmDt_WD1_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_negedge : X01 := '0';
     variable TmDt_WD0_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD5_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD5_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD4_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD4_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD3_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD3_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD2_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD2_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD1_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD1_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD0_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD0_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_negedge : X01 := '0';
     variable TmDt_WEN_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_BLKEN_WCLK_negedge : X01 := '0';
     variable TmDt_BLKEN_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     --type SL_TO_INT is array(std_ulogic range <>) of integer;
     --constant INT :SL_TO_INT('U' to '-') := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;
  
     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable WEN_delayed : std_ulogic := 'X';
     variable REN_delayed : std_ulogic := 'X';
     variable WEN_previous : std_ulogic := 'X';
     variable REN_previous : std_ulogic := 'X';
     variable BLKEN_delayed : std_ulogic := 'X';
     variable BLKEN_previous : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WRAD5_delayed : std_ulogic := 'X';
     variable WRAD4_delayed : std_ulogic := 'X';
     variable WRAD3_delayed : std_ulogic := 'X';
     variable WRAD2_delayed : std_ulogic := 'X';
     variable WRAD1_delayed : std_ulogic := 'X';
     variable WRAD0_delayed : std_ulogic := 'X';
     variable WRAD5_previous : std_ulogic := 'X';
     variable WRAD4_previous : std_ulogic := 'X';
     variable WRAD3_previous : std_ulogic := 'X';
     variable WRAD2_previous : std_ulogic := 'X';
     variable WRAD1_previous : std_ulogic := 'X';
     variable WRAD0_previous : std_ulogic := 'X';
     variable RDAD5_delayed : std_ulogic := 'X';
     variable RDAD4_delayed : std_ulogic := 'X';
     variable RDAD3_delayed : std_ulogic := 'X';
     variable RDAD2_delayed : std_ulogic := 'X';
     variable RDAD1_delayed : std_ulogic := 'X';
     variable RDAD0_delayed : std_ulogic := 'X';
     variable RDAD5_previous : std_ulogic := 'X';
     variable RDAD4_previous : std_ulogic := 'X';
     variable RDAD3_previous : std_ulogic := 'X';
     variable RDAD2_previous : std_ulogic := 'X';
     variable RDAD1_previous : std_ulogic := 'X';
     variable RDAD0_previous : std_ulogic := 'X';
  
  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RDAD high or low before RCLK falling
      --   Hold  RDAD high or low after RCLK falling

      VitalSetupHoldCheck ( Tviol_RDAD5_RCLK_negedge,
                            TmDt_RDAD5_RCLK_negedge,
                            RDAD5_ipd, "RDAD5",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD5_RCLK_noedge_negedge,
                            tsetup_RDAD5_RCLK_noedge_negedge,
                            thold_RDAD5_RCLK_noedge_negedge,
                            thold_RDAD5_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD4_RCLK_negedge,
                            TmDt_RDAD4_RCLK_negedge,
                            RDAD4_ipd, "RDAD4",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD4_RCLK_noedge_negedge,
                            tsetup_RDAD4_RCLK_noedge_negedge,
                            thold_RDAD4_RCLK_noedge_negedge,
                            thold_RDAD4_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD3_RCLK_negedge,
                            TmDt_RDAD3_RCLK_negedge,
                            RDAD3_ipd, "RDAD3",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD3_RCLK_noedge_negedge,
                            tsetup_RDAD3_RCLK_noedge_negedge,
                            thold_RDAD3_RCLK_noedge_negedge,
                            thold_RDAD3_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD2_RCLK_negedge,
                            TmDt_RDAD2_RCLK_negedge,
                            RDAD2_ipd, "RDAD2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD2_RCLK_noedge_negedge,
                            tsetup_RDAD2_RCLK_noedge_negedge,
                            thold_RDAD2_RCLK_noedge_negedge,
                            thold_RDAD2_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD1_RCLK_negedge,
                            TmDt_RDAD1_RCLK_negedge,
                            RDAD1_ipd, "RDAD1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD1_RCLK_noedge_negedge,
                            tsetup_RDAD1_RCLK_noedge_negedge,
                            thold_RDAD1_RCLK_noedge_negedge,
                            thold_RDAD1_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD0_RCLK_negedge,
                            TmDt_RDAD0_RCLK_negedge,
                            RDAD0_ipd, "RDAD0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD0_RCLK_noedge_negedge,
                            tsetup_RDAD0_RCLK_noedge_negedge,
                            thold_RDAD0_RCLK_noedge_negedge,
                            thold_RDAD0_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup REN high before RCLK falling
      --   Hold  REN high after RCLK falling

      VitalSetupHoldCheck ( Tviol_REN_RCLK_negedge,
                            TmDt_REN_RCLK_negedge,
                            REN_ipd, "REN",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_REN_RCLK_noedge_negedge,
                            tsetup_REN_RCLK_noedge_negedge,
                            thold_REN_RCLK_noedge_negedge,
                            thold_REN_RCLK_noedge_negedge,
                            TimingCheckOn,
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup BLKEN high or low before WCLK falling
      --   Hold  BLKEN high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_BLKEN_WCLK_negedge,
                            TmDt_BLKEN_WCLK_negedge,
                            BLKEN_ipd, "BLKEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_BLKEN_WCLK_noedge_negedge,
                            tsetup_BLKEN_WCLK_noedge_negedge,
                            thold_BLKEN_WCLK_noedge_negedge,
                            thold_BLKEN_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WRAD high or low before WCLK falling
      --   Hold  WRAD high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_WRAD5_WCLK_negedge,
                            TmDt_WRAD5_WCLK_negedge,
                            WRAD5_ipd, "WRAD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD5_WCLK_noedge_negedge,
                            tsetup_WRAD5_WCLK_noedge_negedge,
                            thold_WRAD5_WCLK_noedge_negedge,
                            thold_WRAD5_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD4_WCLK_negedge,
                            TmDt_WRAD4_WCLK_negedge,
                            WRAD4_ipd, "WRAD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD4_WCLK_noedge_negedge,
                            tsetup_WRAD4_WCLK_noedge_negedge,
                            thold_WRAD4_WCLK_noedge_negedge,
                            thold_WRAD4_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD3_WCLK_negedge,
                            TmDt_WRAD3_WCLK_negedge,
                            WRAD3_ipd, "WRAD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD3_WCLK_noedge_negedge,
                            tsetup_WRAD3_WCLK_noedge_negedge,
                            thold_WRAD3_WCLK_noedge_negedge,
                            thold_WRAD3_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD2_WCLK_negedge,
                            TmDt_WRAD2_WCLK_negedge,
                            WRAD2_ipd, "WRAD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD2_WCLK_noedge_negedge,
                            tsetup_WRAD2_WCLK_noedge_negedge,
                            thold_WRAD2_WCLK_noedge_negedge,
                            thold_WRAD2_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD1_WCLK_negedge,
                            TmDt_WRAD1_WCLK_negedge,
                            WRAD1_ipd, "WRAD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD1_WCLK_noedge_negedge,
                            tsetup_WRAD1_WCLK_noedge_negedge,
                            thold_WRAD1_WCLK_noedge_negedge,
                            thold_WRAD1_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD0_WCLK_negedge,
                            TmDt_WRAD0_WCLK_negedge,
                            WRAD0_ipd, "WRAD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD0_WCLK_noedge_negedge,
                            tsetup_WRAD0_WCLK_noedge_negedge,
                            thold_WRAD0_WCLK_noedge_negedge,
                            thold_WRAD0_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WD high or low before WCLK falling
      --   Hold  WD high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_negedge,
                            TmDt_WD3_WCLK_negedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_noedge_negedge,
                            tsetup_WD3_WCLK_noedge_negedge,
                            thold_WD3_WCLK_noedge_negedge,
                            thold_WD3_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_negedge,
                            TmDt_WD2_WCLK_negedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_noedge_negedge,
                            tsetup_WD2_WCLK_noedge_negedge,
                            thold_WD2_WCLK_noedge_negedge,
                            thold_WD2_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_negedge,
                            TmDt_WD1_WCLK_negedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_noedge_negedge,
                            tsetup_WD1_WCLK_noedge_negedge,
                            thold_WD1_WCLK_noedge_negedge,
                            thold_WD1_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_negedge,
                            TmDt_WD0_WCLK_negedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_noedge_negedge,
                            tsetup_WD0_WCLK_noedge_negedge,
                            thold_WD0_WCLK_noedge_negedge,
                            thold_WD0_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup WEN high before WCLK falling
      --   Hold  WEN high after WCLK falling

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_negedge,
                            TmDt_WEN_WCLK_negedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_noedge_negedge,
                            tsetup_WEN_WCLK_noedge_negedge,
                            thold_WEN_WCLK_noedge_negedge,
                            thold_WEN_WCLK_noedge_negedge,
                            (To_X01(BLKEN_ipd)=BLKENS),
                            '\',
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM4FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
    
    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      -- Convert Write Address Signal to Integer
      WADDR := ((INT(WRAD5_delayed)*32)+(INT(WRAD4_delayed)*16)+(INT(WRAD3_delayed)*8)+
		(INT(WRAD2_delayed)*4)+(INT(WRAD1_delayed)*2)+(INT(WRAD0_delayed)));

      if (TO_X01(WCLK_ipd)='X') then
        if (TO_X01(WCLK_previous) /= 'X') then
	  assert false
	  report ": WCLK unknown"
	  severity Warning;
	end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='0')) then
	case TO_X01(WEN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (TO_X01(BLKEN_delayed) = 'X') then
              if (TO_X01(BLKEN_previous) /= 'X') then
	        assert false
	        report ": BLKEN unknown"
	        severity Warning;
	      end if;
	    elsif (TO_X01(BLKEN_delayed) = BLKENS) then
	      if (WADDR < 0) then
		if (TO_X01(WRAD5_delayed) = 'X') and (TO_X01(WRAD5_previous) /= 'X') then
		  assert false
		  report ": WRAD5 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD4_delayed) = 'X') and (TO_X01(WRAD4_previous) /= 'X') then
		  assert false
		  report ": WRAD4 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD3_delayed) = 'X') and (TO_X01(WRAD3_previous) /= 'X') then
		  assert false
		  report ": WRAD3 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD2_delayed) = 'X') and (TO_X01(WRAD2_previous) /= 'X') then
		  assert false
		  report ": WRAD2 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD1_delayed) = 'X') and (TO_X01(WRAD1_previous) /= 'X') then
		  assert false
		  report ": WRAD1 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD0_delayed) = 'X') and (TO_X01(WRAD0_previous) /= 'X') then
		  assert false
		  report ": WRAD0 unknown"
		  severity Warning;
		end if;
	      else 
		RAM_TMP(WADDR) <= WD3_delayed & WD2_delayed & WD1_delayed & WD0_delayed ; 
	      end if;
	    else
	      null;
	    end if;
	  when others =>
            if (TO_X01(WEN_previous) /= 'X') then
	      assert false
	      report ": WEN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      -- Convert Read Address Signal to Integer
      RADDR := ((INT(RDAD5_delayed)*32)+(INT(RDAD4_delayed)*16)+(INT(RDAD3_delayed)*8)+
		(INT(RDAD2_delayed)*4)+(INT(RDAD1_delayed)*2)+(INT(RDAD0_delayed)));

      if (TO_X01(RCLK_ipd) = 'X') then
	RD3_zd := 'X';
	RD2_zd := 'X';
	RD1_zd := 'X';
	RD0_zd := 'X';
	if (TO_X01(RCLK_previous) /= 'X') then
	  assert false
	  report ": RCLK unknown"
	  severity Warning;
	end if;
      elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '0')) then
	case TO_X01(REN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (RADDR < 0) then
	      RD3_zd := 'X';
	      RD2_zd := 'X';
	      RD1_zd := 'X';
	      RD0_zd := 'X';
	      if (TO_X01(RDAD5_delayed) = 'X') and (TO_X01(RDAD5_previous) /= 'X') then
		assert false
		report ": RDAD5 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD4_delayed) = 'X') and (TO_X01(RDAD4_previous) /= 'X') then
		assert false
		report ": RDAD4 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD3_delayed) = 'X') and (TO_X01(RDAD3_previous) /= 'X') then
		assert false
		report ": RDAD3 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD2_delayed) = 'X') and (TO_X01(RDAD2_previous) /= 'X') then
		assert false
		report ": RDAD2 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD1_delayed) = 'X') and (TO_X01(RDAD1_previous) /= 'X') then
		assert false
		report ": RDAD1 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD0_delayed) = 'X') and (TO_X01(RDAD0_previous) /= 'X') then
		assert false
		report ": RDAD0 unknown"
		severity Warning;
	      end if;
	    else
	      RD3_zd := RAM_TMP(RADDR)(3);
	      RD2_zd := RAM_TMP(RADDR)(2);
	      RD1_zd := RAM_TMP(RADDR)(1);
	      RD0_zd := RAM_TMP(RADDR)(0);
	    end if;
	  when others =>
	    RD3_zd := 'X';
	    RD2_zd := 'X';
	    RD1_zd := 'X';
	    RD0_zd := 'X';
            if (TO_X01(REN_previous) /= 'X') then
	      assert false
	      report ": REN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;
      
      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      WEN_previous := WEN_delayed;
      REN_previous := REN_delayed;
      WEN_delayed := WEN_ipd;
      REN_delayed := REN_ipd;
      BLKEN_previous := BLKEN_delayed;
      BLKEN_delayed := BLKEN_ipd;
      WD3_delayed := WD3_ipd;
      WD2_delayed := WD2_ipd;
      WD1_delayed := WD1_ipd;
      WD0_delayed := WD0_ipd;
      WRAD5_previous := WRAD5_delayed;
      WRAD4_previous := WRAD4_delayed;
      WRAD3_previous := WRAD3_delayed;
      WRAD2_previous := WRAD2_delayed;
      WRAD1_previous := WRAD1_delayed;
      WRAD0_previous := WRAD0_delayed;
      WRAD5_delayed := WRAD5_ipd;
      WRAD4_delayed := WRAD4_ipd;
      WRAD3_delayed := WRAD3_ipd;
      WRAD2_delayed := WRAD2_ipd;
      WRAD1_delayed := WRAD1_ipd;
      WRAD0_delayed := WRAD0_ipd;
      RDAD5_previous := RDAD5_delayed;
      RDAD4_previous := RDAD4_delayed;
      RDAD3_previous := RDAD3_delayed;
      RDAD2_previous := RDAD2_delayed;
      RDAD1_previous := RDAD1_delayed;
      RDAD0_previous := RDAD0_delayed;
      RDAD5_delayed := RDAD5_ipd;
      RDAD4_delayed := RDAD4_ipd;
      RDAD3_delayed := RDAD3_ipd;
      RDAD2_delayed := RDAD2_ipd;
      RDAD1_delayed := RDAD1_ipd;
      RDAD0_delayed := RDAD0_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD3,
	GlitchData => RD3_GlitchData,
	OutSignalName => "RD3",
	OutTemp => RD3_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD3), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD2,
	GlitchData => RD2_GlitchData,
	OutSignalName => "RD2",
	OutTemp => RD2_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD2), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD1,
	GlitchData => RD1_GlitchData,
	OutSignalName => "RD1",
	OutTemp => RD1_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD1), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD0,
	GlitchData => RD0_GlitchData,
	OutSignalName => "RD0",
	OutTemp => RD0_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD0), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

  end process VITALBehavior;

end VITAL_ACT;
-----------------------------------------------------------------
--  Proxy Modeling, Inc. 
--
--  Actel RAM4FR VHDL behavioral model
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - Jan/22/96 - Initial Delivery
-- 1.1 - 12/6/96 by DNW - Modified SL_TO_INT.
-- 1.2 - 3/3/97 by DNW - WDx_delayed variables added.
-- 1.3 - 3/6/98 by DNW - Issue "unknown" msg. only if 0/1->X Xtion.
-- 1.4 - 5/27/98 by DNW - Initaialize _ipd signals to X instead of 0.
-- 
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity RAM4FR is
  GENERIC (
        tipd_RDAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD5_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of RAM4FR : entity is TRUE;
  
end RAM4FR;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM4FR is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal WRAD5_ipd : std_ulogic := 'X';
  signal WRAD4_ipd : std_ulogic := 'X';
  signal WRAD3_ipd : std_ulogic := 'X';
  signal WRAD2_ipd : std_ulogic := 'X';
  signal WRAD1_ipd : std_ulogic := 'X';
  signal WRAD0_ipd : std_ulogic := 'X';
  signal WD3_ipd : std_ulogic := 'X';
  signal WD2_ipd : std_ulogic := 'X';
  signal WD1_ipd : std_ulogic := 'X';
  signal WD0_ipd : std_ulogic := 'X';
  signal RDAD5_ipd : std_ulogic := 'X';
  signal RDAD4_ipd : std_ulogic := 'X';
  signal RDAD3_ipd : std_ulogic := 'X';
  signal RDAD2_ipd : std_ulogic := 'X';
  signal RDAD1_ipd : std_ulogic := 'X';
  signal RDAD0_ipd : std_ulogic := 'X';
  signal BLKEN_ipd : std_ulogic := 'X';
  signal WEN_ipd : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal REN_ipd : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  type MEM is array(0 to 63) of std_ulogic_vector(3 downto 0);
   signal RAM_TMP : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (WRAD5_ipd, WRAD5, VitalExtendToFillDelay(tipd_WRAD5));
    VitalWireDelay (WRAD4_ipd, WRAD4, VitalExtendToFillDelay(tipd_WRAD4));
    VitalWireDelay (WRAD3_ipd, WRAD3, VitalExtendToFillDelay(tipd_WRAD3));
    VitalWireDelay (WRAD2_ipd, WRAD2, VitalExtendToFillDelay(tipd_WRAD2));
    VitalWireDelay (WRAD1_ipd, WRAD1, VitalExtendToFillDelay(tipd_WRAD1));
    VitalWireDelay (WRAD0_ipd, WRAD0, VitalExtendToFillDelay(tipd_WRAD0));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (RDAD5_ipd, RDAD5, VitalExtendToFillDelay(tipd_RDAD5));
    VitalWireDelay (RDAD4_ipd, RDAD4, VitalExtendToFillDelay(tipd_RDAD4));
    VitalWireDelay (RDAD3_ipd, RDAD3, VitalExtendToFillDelay(tipd_RDAD3));
    VitalWireDelay (RDAD2_ipd, RDAD2, VitalExtendToFillDelay(tipd_RDAD2));
    VitalWireDelay (RDAD1_ipd, RDAD1, VitalExtendToFillDelay(tipd_RDAD1));
    VitalWireDelay (RDAD0_ipd, RDAD0, VitalExtendToFillDelay(tipd_RDAD0));
    VitalWireDelay (BLKEN_ipd, BLKEN, VitalExtendToFillDelay(tipd_BLKEN));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (REN_ipd, REN, VitalExtendToFillDelay(tipd_REN));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (RDAD5_ipd, RDAD4_ipd, RDAD3_ipd, RDAD2_ipd, 
		RDAD1_ipd, RDAD0_ipd, REN_ipd, RCLK_ipd, 
		WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd, WRAD5_ipd, WRAD4_ipd, 
		WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, WEN_ipd, 
		BLKEN_ipd, BLKENS, WCLK_ipd)

     --  Read Timing Check Results
     variable Tviol_RDAD5_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD5_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD4_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD4_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD3_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD2_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD1_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD0_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_REN_RCLK_posedge : X01 := '0';
     variable TmDt_REN_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_WD3_WCLK_negedge : X01 := '0';
     variable TmDt_WD3_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_negedge : X01 := '0';
     variable TmDt_WD2_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_negedge : X01 := '0';
     variable TmDt_WD1_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_negedge : X01 := '0';
     variable TmDt_WD0_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD5_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD5_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD4_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD4_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD3_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD3_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD2_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD2_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD1_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD1_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD0_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD0_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_negedge : X01 := '0';
     variable TmDt_WEN_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_BLKEN_WCLK_negedge : X01 := '0';
     variable TmDt_BLKEN_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     --type SL_TO_INT is array(std_ulogic range <>) of integer;
     --constant INT :SL_TO_INT('U' to '-') := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;
  
     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable WEN_delayed : std_ulogic := 'X';
     variable REN_delayed : std_ulogic := 'X';
     variable WEN_previous : std_ulogic := 'X';
     variable REN_previous : std_ulogic := 'X';
     variable BLKEN_delayed : std_ulogic := 'X';
     variable BLKEN_previous : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WRAD5_delayed : std_ulogic := 'X';
     variable WRAD4_delayed : std_ulogic := 'X';
     variable WRAD3_delayed : std_ulogic := 'X';
     variable WRAD2_delayed : std_ulogic := 'X';
     variable WRAD1_delayed : std_ulogic := 'X';
     variable WRAD0_delayed : std_ulogic := 'X';
     variable WRAD5_previous : std_ulogic := 'X';
     variable WRAD4_previous : std_ulogic := 'X';
     variable WRAD3_previous : std_ulogic := 'X';
     variable WRAD2_previous : std_ulogic := 'X';
     variable WRAD1_previous : std_ulogic := 'X';
     variable WRAD0_previous : std_ulogic := 'X';
     variable RDAD5_delayed : std_ulogic := 'X';
     variable RDAD4_delayed : std_ulogic := 'X';
     variable RDAD3_delayed : std_ulogic := 'X';
     variable RDAD2_delayed : std_ulogic := 'X';
     variable RDAD1_delayed : std_ulogic := 'X';
     variable RDAD0_delayed : std_ulogic := 'X';
     variable RDAD5_previous : std_ulogic := 'X';
     variable RDAD4_previous : std_ulogic := 'X';
     variable RDAD3_previous : std_ulogic := 'X';
     variable RDAD2_previous : std_ulogic := 'X';
     variable RDAD1_previous : std_ulogic := 'X';
     variable RDAD0_previous : std_ulogic := 'X';
  
  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RDAD high or low before RCLK rising
      --   Hold  RDAD high or low after RCLK rising

      VitalSetupHoldCheck ( Tviol_RDAD5_RCLK_posedge,
                            TmDt_RDAD5_RCLK_posedge,
                            RDAD5_ipd, "RDAD5",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD5_RCLK_noedge_posedge,
                            tsetup_RDAD5_RCLK_noedge_posedge,
                            thold_RDAD5_RCLK_noedge_posedge,
                            thold_RDAD5_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD4_RCLK_posedge,
                            TmDt_RDAD4_RCLK_posedge,
                            RDAD4_ipd, "RDAD4",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD4_RCLK_noedge_posedge,
                            tsetup_RDAD4_RCLK_noedge_posedge,
                            thold_RDAD4_RCLK_noedge_posedge,
                            thold_RDAD4_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD3_RCLK_posedge,
                            TmDt_RDAD3_RCLK_posedge,
                            RDAD3_ipd, "RDAD3",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD3_RCLK_noedge_posedge,
                            tsetup_RDAD3_RCLK_noedge_posedge,
                            thold_RDAD3_RCLK_noedge_posedge,
                            thold_RDAD3_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD2_RCLK_posedge,
                            TmDt_RDAD2_RCLK_posedge,
                            RDAD2_ipd, "RDAD2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD2_RCLK_noedge_posedge,
                            tsetup_RDAD2_RCLK_noedge_posedge,
                            thold_RDAD2_RCLK_noedge_posedge,
                            thold_RDAD2_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD1_RCLK_posedge,
                            TmDt_RDAD1_RCLK_posedge,
                            RDAD1_ipd, "RDAD1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD1_RCLK_noedge_posedge,
                            tsetup_RDAD1_RCLK_noedge_posedge,
                            thold_RDAD1_RCLK_noedge_posedge,
                            thold_RDAD1_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD0_RCLK_posedge,
                            TmDt_RDAD0_RCLK_posedge,
                            RDAD0_ipd, "RDAD0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD0_RCLK_noedge_posedge,
                            tsetup_RDAD0_RCLK_noedge_posedge,
                            thold_RDAD0_RCLK_noedge_posedge,
                            thold_RDAD0_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup REN high before RCLK rising
      --   Hold  REN high after RCLK rising

      VitalSetupHoldCheck ( Tviol_REN_RCLK_posedge,
                            TmDt_REN_RCLK_posedge,
                            REN_ipd, "REN",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_REN_RCLK_noedge_posedge,
                            tsetup_REN_RCLK_noedge_posedge,
                            thold_REN_RCLK_noedge_posedge,
                            thold_REN_RCLK_noedge_posedge,
                            TimingCheckOn,
                            '/',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup BLKEN high or low before WCLK falling
      --   Hold  BLKEN high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_BLKEN_WCLK_negedge,
                            TmDt_BLKEN_WCLK_negedge,
                            BLKEN_ipd, "BLKEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_BLKEN_WCLK_noedge_negedge,
                            tsetup_BLKEN_WCLK_noedge_negedge,
                            thold_BLKEN_WCLK_noedge_negedge,
                            thold_BLKEN_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WRAD high or low before WCLK falling
      --   Hold  WRAD high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_WRAD5_WCLK_negedge,
                            TmDt_WRAD5_WCLK_negedge,
                            WRAD5_ipd, "WRAD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD5_WCLK_noedge_negedge,
                            tsetup_WRAD5_WCLK_noedge_negedge,
                            thold_WRAD5_WCLK_noedge_negedge,
                            thold_WRAD5_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD4_WCLK_negedge,
                            TmDt_WRAD4_WCLK_negedge,
                            WRAD4_ipd, "WRAD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD4_WCLK_noedge_negedge,
                            tsetup_WRAD4_WCLK_noedge_negedge,
                            thold_WRAD4_WCLK_noedge_negedge,
                            thold_WRAD4_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD3_WCLK_negedge,
                            TmDt_WRAD3_WCLK_negedge,
                            WRAD3_ipd, "WRAD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD3_WCLK_noedge_negedge,
                            tsetup_WRAD3_WCLK_noedge_negedge,
                            thold_WRAD3_WCLK_noedge_negedge,
                            thold_WRAD3_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD2_WCLK_negedge,
                            TmDt_WRAD2_WCLK_negedge,
                            WRAD2_ipd, "WRAD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD2_WCLK_noedge_negedge,
                            tsetup_WRAD2_WCLK_noedge_negedge,
                            thold_WRAD2_WCLK_noedge_negedge,
                            thold_WRAD2_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD1_WCLK_negedge,
                            TmDt_WRAD1_WCLK_negedge,
                            WRAD1_ipd, "WRAD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD1_WCLK_noedge_negedge,
                            tsetup_WRAD1_WCLK_noedge_negedge,
                            thold_WRAD1_WCLK_noedge_negedge,
                            thold_WRAD1_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD0_WCLK_negedge,
                            TmDt_WRAD0_WCLK_negedge,
                            WRAD0_ipd, "WRAD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD0_WCLK_noedge_negedge,
                            tsetup_WRAD0_WCLK_noedge_negedge,
                            thold_WRAD0_WCLK_noedge_negedge,
                            thold_WRAD0_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WD high or low before WCLK falling
      --   Hold  WD high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_negedge,
                            TmDt_WD3_WCLK_negedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_noedge_negedge,
                            tsetup_WD3_WCLK_noedge_negedge,
                            thold_WD3_WCLK_noedge_negedge,
                            thold_WD3_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_negedge,
                            TmDt_WD2_WCLK_negedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_noedge_negedge,
                            tsetup_WD2_WCLK_noedge_negedge,
                            thold_WD2_WCLK_noedge_negedge,
                            thold_WD2_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_negedge,
                            TmDt_WD1_WCLK_negedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_noedge_negedge,
                            tsetup_WD1_WCLK_noedge_negedge,
                            thold_WD1_WCLK_noedge_negedge,
                            thold_WD1_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_negedge,
                            TmDt_WD0_WCLK_negedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_noedge_negedge,
                            tsetup_WD0_WCLK_noedge_negedge,
                            thold_WD0_WCLK_noedge_negedge,
                            thold_WD0_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup WEN high before WCLK falling
      --   Hold  WEN high after WCLK falling

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_negedge,
                            TmDt_WEN_WCLK_negedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_noedge_negedge,
                            tsetup_WEN_WCLK_noedge_negedge,
                            thold_WEN_WCLK_noedge_negedge,
                            thold_WEN_WCLK_noedge_negedge,
                            TimingCheckOn,
                            '\',
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM4FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
    
    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      -- Convert Write Address Signal to Integer
      WADDR := ((INT(WRAD5_delayed)*32)+(INT(WRAD4_delayed)*16)+(INT(WRAD3_delayed)*8)+
		(INT(WRAD2_delayed)*4)+(INT(WRAD1_delayed)*2)+(INT(WRAD0_delayed)));

      if (TO_X01(WCLK_ipd)='X') then
        if (TO_X01(WCLK_previous) /= 'X') then
	  assert false
	  report ": WCLK unknown"
	  severity Warning;
	end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='0')) then
	case TO_X01(WEN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (TO_X01(BLKEN_delayed) = 'X') then
              if (TO_X01(BLKEN_previous) /= 'X') then
	        assert false
	        report ": BLKEN unknown"
	        severity Warning;
	      end if;
	    elsif (TO_X01(BLKEN_delayed) = BLKENS) then
	      if (WADDR < 0) then
		if (TO_X01(WRAD5_delayed) = 'X') and (TO_X01(WRAD5_previous) /= 'X') then
		  assert false
		  report ": WRAD5 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD4_delayed) = 'X') and (TO_X01(WRAD4_previous) /= 'X') then
		  assert false
		  report ": WRAD4 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD3_delayed) = 'X') and (TO_X01(WRAD3_previous) /= 'X') then
		  assert false
		  report ": WRAD3 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD2_delayed) = 'X') and (TO_X01(WRAD2_previous) /= 'X') then
		  assert false
		  report ": WRAD2 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD1_delayed) = 'X') and (TO_X01(WRAD1_previous) /= 'X') then
		  assert false
		  report ": WRAD1 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD0_delayed) = 'X') and (TO_X01(WRAD0_previous) /= 'X') then
		  assert false
		  report ": WRAD0 unknown"
		  severity Warning;
		end if;
	      else 
		RAM_TMP(WADDR) <= WD3_delayed & WD2_delayed & WD1_delayed & WD0_delayed ; 
	      end if;
	    else
	      null;
	    end if;
	  when others =>
            if (TO_X01(WEN_previous) /= 'X') then
	      assert false
	      report ": WEN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      -- Convert Read Address Signal to Integer
      RADDR := ((INT(RDAD5_delayed)*32)+(INT(RDAD4_delayed)*16)+(INT(RDAD3_delayed)*8)+
		(INT(RDAD2_delayed)*4)+(INT(RDAD1_delayed)*2)+(INT(RDAD0_delayed)));

      if (TO_X01(RCLK_ipd) = 'X') then
	RD3_zd := 'X';
	RD2_zd := 'X';
	RD1_zd := 'X';
	RD0_zd := 'X';
	if (TO_X01(RCLK_previous) /= 'X') then
	  assert false
	  report ": RCLK unknown"
	  severity Warning;
	end if;
      elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1')) then
	case TO_X01(REN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (RADDR < 0) then
	      RD3_zd := 'X';
	      RD2_zd := 'X';
	      RD1_zd := 'X';
	      RD0_zd := 'X';
	      if (TO_X01(RDAD5_delayed) = 'X') and (TO_X01(RDAD5_previous) /= 'X') then
		assert false
		report ": RDAD5 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD4_delayed) = 'X') and (TO_X01(RDAD4_previous) /= 'X') then
		assert false
		report ": RDAD4 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD3_delayed) = 'X') and (TO_X01(RDAD3_previous) /= 'X') then
		assert false
		report ": RDAD3 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD2_delayed) = 'X') and (TO_X01(RDAD2_previous) /= 'X') then
		assert false
		report ": RDAD2 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD1_delayed) = 'X') and (TO_X01(RDAD1_previous) /= 'X') then
		assert false
		report ": RDAD1 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD0_delayed) = 'X') and (TO_X01(RDAD0_previous) /= 'X') then
		assert false
		report ": RDAD0 unknown"
		severity Warning;
	      end if;
	    else
	      RD3_zd := RAM_TMP(RADDR)(3);
	      RD2_zd := RAM_TMP(RADDR)(2);
	      RD1_zd := RAM_TMP(RADDR)(1);
	      RD0_zd := RAM_TMP(RADDR)(0);
	    end if;
	  when others =>
	    RD3_zd := 'X';
	    RD2_zd := 'X';
	    RD1_zd := 'X';
	    RD0_zd := 'X';
            if (TO_X01(REN_previous) /= 'X') then
	      assert false
	      report ": REN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;
      
      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      WEN_previous := WEN_delayed;
      REN_previous := REN_delayed;
      WEN_delayed := WEN_ipd;
      REN_delayed := REN_ipd;
      BLKEN_previous := BLKEN_delayed;
      BLKEN_delayed := BLKEN_ipd;
      WD3_delayed := WD3_ipd;
      WD2_delayed := WD2_ipd;
      WD1_delayed := WD1_ipd;
      WD0_delayed := WD0_ipd;
      WRAD5_previous := WRAD5_delayed;
      WRAD4_previous := WRAD4_delayed;
      WRAD3_previous := WRAD3_delayed;
      WRAD2_previous := WRAD2_delayed;
      WRAD1_previous := WRAD1_delayed;
      WRAD0_previous := WRAD0_delayed;
      WRAD5_delayed := WRAD5_ipd;
      WRAD4_delayed := WRAD4_ipd;
      WRAD3_delayed := WRAD3_ipd;
      WRAD2_delayed := WRAD2_ipd;
      WRAD1_delayed := WRAD1_ipd;
      WRAD0_delayed := WRAD0_ipd;
      RDAD5_previous := RDAD5_delayed;
      RDAD4_previous := RDAD4_delayed;
      RDAD3_previous := RDAD3_delayed;
      RDAD2_previous := RDAD2_delayed;
      RDAD1_previous := RDAD1_delayed;
      RDAD0_previous := RDAD0_delayed;
      RDAD5_delayed := RDAD5_ipd;
      RDAD4_delayed := RDAD4_ipd;
      RDAD3_delayed := RDAD3_ipd;
      RDAD2_delayed := RDAD2_ipd;
      RDAD1_delayed := RDAD1_ipd;
      RDAD0_delayed := RDAD0_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD3,
	GlitchData => RD3_GlitchData,
	OutSignalName => "RD3",
	OutTemp => RD3_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD3), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD2,
	GlitchData => RD2_GlitchData,
	OutSignalName => "RD2",
	OutTemp => RD2_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD2), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD1,
	GlitchData => RD1_GlitchData,
	OutSignalName => "RD1",
	OutTemp => RD1_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD1), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD0,
	GlitchData => RD0_GlitchData,
	OutSignalName => "RD0",
	OutTemp => RD0_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD0), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

  end process VITALBehavior;

end VITAL_ACT;
-----------------------------------------------------------------
--  Proxy Modeling, Inc. 
--
--  Actel RAM4RA VHDL behavioral model
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - Jan/22/96 - Initial Delivery
-- 1.1 - 12/6/96 by DNW - Modified SL_TO_INT.
-- 1.2 - 3/3/97 by DNW - WDx_delayed variables added.
-- 1.3 - 3/6/98 by DNW - Issue "unknown" msg. only if 0/1->X Xtion.
-- 1.4 - 5/27/98 by DNW - Initaialize _ipd signals to X instead of 0.
-- 
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity RAM4RA is
  GENERIC (
        tipd_RDAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RDAD5_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD5_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD5_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD5_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_WRAD5_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of RAM4RA : entity is TRUE;
  
end RAM4RA;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM4RA is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal WRAD5_ipd : std_ulogic := 'X';
  signal WRAD4_ipd : std_ulogic := 'X';
  signal WRAD3_ipd : std_ulogic := 'X';
  signal WRAD2_ipd : std_ulogic := 'X';
  signal WRAD1_ipd : std_ulogic := 'X';
  signal WRAD0_ipd : std_ulogic := 'X';
  signal WD3_ipd : std_ulogic := 'X';
  signal WD2_ipd : std_ulogic := 'X';
  signal WD1_ipd : std_ulogic := 'X';
  signal WD0_ipd : std_ulogic := 'X';
  signal RDAD5_ipd : std_ulogic := 'X';
  signal RDAD4_ipd : std_ulogic := 'X';
  signal RDAD3_ipd : std_ulogic := 'X';
  signal RDAD2_ipd : std_ulogic := 'X';
  signal RDAD1_ipd : std_ulogic := 'X';
  signal RDAD0_ipd : std_ulogic := 'X';
  signal BLKEN_ipd : std_ulogic := 'X';
  signal WEN_ipd : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  type MEM is array(0 to 63) of std_ulogic_vector(3 downto 0);
   signal RAM_TMP : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (WRAD5_ipd, WRAD5, VitalExtendToFillDelay(tipd_WRAD5));
    VitalWireDelay (WRAD4_ipd, WRAD4, VitalExtendToFillDelay(tipd_WRAD4));
    VitalWireDelay (WRAD3_ipd, WRAD3, VitalExtendToFillDelay(tipd_WRAD3));
    VitalWireDelay (WRAD2_ipd, WRAD2, VitalExtendToFillDelay(tipd_WRAD2));
    VitalWireDelay (WRAD1_ipd, WRAD1, VitalExtendToFillDelay(tipd_WRAD1));
    VitalWireDelay (WRAD0_ipd, WRAD0, VitalExtendToFillDelay(tipd_WRAD0));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (RDAD5_ipd, RDAD5, VitalExtendToFillDelay(tipd_RDAD5));
    VitalWireDelay (RDAD4_ipd, RDAD4, VitalExtendToFillDelay(tipd_RDAD4));
    VitalWireDelay (RDAD3_ipd, RDAD3, VitalExtendToFillDelay(tipd_RDAD3));
    VitalWireDelay (RDAD2_ipd, RDAD2, VitalExtendToFillDelay(tipd_RDAD2));
    VitalWireDelay (RDAD1_ipd, RDAD1, VitalExtendToFillDelay(tipd_RDAD1));
    VitalWireDelay (RDAD0_ipd, RDAD0, VitalExtendToFillDelay(tipd_RDAD0));
    VitalWireDelay (BLKEN_ipd, BLKEN, VitalExtendToFillDelay(tipd_BLKEN));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (RDAD5_ipd, RDAD4_ipd, RDAD3_ipd, RDAD2_ipd, 
		RDAD1_ipd, RDAD0_ipd, 
		WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd, WRAD5_ipd, WRAD4_ipd, 
		WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, WEN_ipd, 
		BLKEN_ipd, BLKENS, WCLK_ipd, RAM_TMP)

     --  Write Timing Check Results
     variable Tviol_WD3_WCLK_posedge : X01 := '0';
     variable TmDT_WD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_posedge : X01 := '0';
     variable TmDT_WD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_posedge : X01 := '0';
     variable TmDT_WD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_posedge : X01 := '0';
     variable TmDT_WD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD5_WCLK_posedge : X01 := '0';
     variable TmDT_WRAD5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD4_WCLK_posedge : X01 := '0';
     variable TmDT_WRAD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD3_WCLK_posedge : X01 := '0';
     variable TmDT_WRAD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD2_WCLK_posedge : X01 := '0';
     variable TmDT_WRAD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD1_WCLK_posedge : X01 := '0';
     variable TmDT_WRAD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD0_WCLK_posedge : X01 := '0';
     variable TmDT_WRAD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_posedge : X01 := '0';
     variable TmDT_WEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_BLKEN_WCLK_posedge : X01 := '0';
     variable TmDT_BLKEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     --type SL_TO_INT is array(std_ulogic range <>) of integer;
     --constant INT :SL_TO_INT('U' to '-') := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;
  
     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable WEN_delayed : std_ulogic := 'X';
     variable WEN_previous : std_ulogic := 'X';
     variable BLKEN_delayed : std_ulogic := 'X';
     variable BLKEN_previous : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WRAD5_delayed : std_ulogic := 'X';
     variable WRAD4_delayed : std_ulogic := 'X';
     variable WRAD3_delayed : std_ulogic := 'X';
     variable WRAD2_delayed : std_ulogic := 'X';
     variable WRAD1_delayed : std_ulogic := 'X';
     variable WRAD0_delayed : std_ulogic := 'X';
     variable WRAD5_previous : std_ulogic := 'X';
     variable WRAD4_previous : std_ulogic := 'X';
     variable WRAD3_previous : std_ulogic := 'X';
     variable WRAD2_previous : std_ulogic := 'X';
     variable WRAD1_previous : std_ulogic := 'X';
     variable WRAD0_previous : std_ulogic := 'X';
     variable RDAD5_previous : std_ulogic := 'X';
     variable RDAD4_previous : std_ulogic := 'X';
     variable RDAD3_previous : std_ulogic := 'X';
     variable RDAD2_previous : std_ulogic := 'X';
     variable RDAD1_previous : std_ulogic := 'X';
     variable RDAD0_previous : std_ulogic := 'X';
  
  begin  --  process VITALBehavior 

    if (TimingCheckOn) then

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup BLKEN high or low before WCLK rising
      --   Hold  BLKEN high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_BLKEN_WCLK_posedge,
                            TmDT_BLKEN_WCLK_posedge,
                            BLKEN_ipd, "BLKEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_BLKEN_WCLK_noedge_posedge,
                            tsetup_BLKEN_WCLK_noedge_posedge,
                            thold_BLKEN_WCLK_noedge_posedge,
                            thold_BLKEN_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WRAD high or low before WCLK rising
      --   Hold  WRAD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WRAD5_WCLK_posedge,
                            TmDT_WRAD5_WCLK_posedge,
                            WRAD5_ipd, "WRAD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD5_WCLK_noedge_posedge,
                            tsetup_WRAD5_WCLK_noedge_posedge,
                            thold_WRAD5_WCLK_noedge_posedge,
                            thold_WRAD5_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD4_WCLK_posedge,
                            TmDT_WRAD4_WCLK_posedge,
                            WRAD4_ipd, "WRAD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD4_WCLK_noedge_posedge,
                            tsetup_WRAD4_WCLK_noedge_posedge,
                            thold_WRAD4_WCLK_noedge_posedge,
                            thold_WRAD4_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD3_WCLK_posedge,
                            TmDT_WRAD3_WCLK_posedge,
                            WRAD3_ipd, "WRAD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD3_WCLK_noedge_posedge,
                            tsetup_WRAD3_WCLK_noedge_posedge,
                            thold_WRAD3_WCLK_noedge_posedge,
                            thold_WRAD3_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD2_WCLK_posedge,
                            TmDT_WRAD2_WCLK_posedge,
                            WRAD2_ipd, "WRAD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD2_WCLK_noedge_posedge,
                            tsetup_WRAD2_WCLK_noedge_posedge,
                            thold_WRAD2_WCLK_noedge_posedge,
                            thold_WRAD2_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD1_WCLK_posedge,
                            TmDT_WRAD1_WCLK_posedge,
                            WRAD1_ipd, "WRAD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD1_WCLK_noedge_posedge,
                            tsetup_WRAD1_WCLK_noedge_posedge,
                            thold_WRAD1_WCLK_noedge_posedge,
                            thold_WRAD1_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD0_WCLK_posedge,
                            TmDT_WRAD0_WCLK_posedge,
                            WRAD0_ipd, "WRAD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD0_WCLK_noedge_posedge,
                            tsetup_WRAD0_WCLK_noedge_posedge,
                            thold_WRAD0_WCLK_noedge_posedge,
                            thold_WRAD0_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WD high or low before WCLK rising
      --   Hold  WD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_posedge,
                            TmDT_WD3_WCLK_posedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_noedge_posedge,
                            tsetup_WD3_WCLK_noedge_posedge,
                            thold_WD3_WCLK_noedge_posedge,
                            thold_WD3_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_posedge,
                            TmDT_WD2_WCLK_posedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_noedge_posedge,
                            tsetup_WD2_WCLK_noedge_posedge,
                            thold_WD2_WCLK_noedge_posedge,
                            thold_WD2_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_posedge,
                            TmDT_WD1_WCLK_posedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_noedge_posedge,
                            tsetup_WD1_WCLK_noedge_posedge,
                            thold_WD1_WCLK_noedge_posedge,
                            thold_WD1_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_posedge,
                            TmDT_WD0_WCLK_posedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_noedge_posedge,
                            tsetup_WD0_WCLK_noedge_posedge,
                            thold_WD0_WCLK_noedge_posedge,
                            thold_WD0_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup WEN high before WCLK rising
      --   Hold  WEN high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_posedge,
                            TmDT_WEN_WCLK_posedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_noedge_posedge,
                            tsetup_WEN_WCLK_noedge_posedge,
                            thold_WEN_WCLK_noedge_posedge,
                            thold_WEN_WCLK_noedge_posedge,
                            (To_X01(BLKEN_ipd)=BLKENS),
                            '/',
                            InstancePath & "/RAM4RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM4RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
    
    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      -- Convert Write Address Signal to Integer
      WADDR := ((INT(WRAD5_delayed)*32)+(INT(WRAD4_delayed)*16)+(INT(WRAD3_delayed)*8)+
		(INT(WRAD2_delayed)*4)+(INT(WRAD1_delayed)*2)+(INT(WRAD0_delayed)));

      if (TO_X01(WCLK_ipd)='X') then
        if (TO_X01(WCLK_previous) /= 'X') then
	  assert false
	  report ": WCLK unknown"
	  severity Warning;
	end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	case TO_X01(WEN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (TO_X01(BLKEN_delayed) = 'X') then
              if (TO_X01(BLKEN_previous) /= 'X') then
	        assert false
	        report ": BLKEN unknown"
	        severity Warning;
	      end if;
	    elsif (TO_X01(BLKEN_delayed) = BLKENS) then
	      if (WADDR < 0) then
		if (TO_X01(WRAD5_delayed) = 'X') and (TO_X01(WRAD5_previous) /= 'X') then
		  assert false
		  report ": WRAD5 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD4_delayed) = 'X') and (TO_X01(WRAD4_previous) /= 'X') then
		  assert false
		  report ": WRAD4 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD3_delayed) = 'X') and (TO_X01(WRAD3_previous) /= 'X') then
		  assert false
		  report ": WRAD3 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD2_delayed) = 'X') and (TO_X01(WRAD2_previous) /= 'X') then
		  assert false
		  report ": WRAD2 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD1_delayed) = 'X') and (TO_X01(WRAD1_previous) /= 'X') then
		  assert false
		  report ": WRAD1 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD0_delayed) = 'X') and (TO_X01(WRAD0_previous) /= 'X') then
		  assert false
		  report ": WRAD0 unknown"
		  severity Warning;
		end if;
	      else 
		RAM_TMP(WADDR) <= WD3_delayed & WD2_delayed & WD1_delayed & WD0_delayed ; 
	      end if;
	    else
	      null;
	    end if;
	  when others =>
            if (TO_X01(WEN_previous) /= 'X') then
	      assert false
	      report ": WEN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      -- Convert Read Address Signal to Integer
      RADDR := ((INT(RDAD5_ipd)*32)+(INT(RDAD4_ipd)*16)+(INT(RDAD3_ipd)*8)+
		(INT(RDAD2_ipd)*4)+(INT(RDAD1_ipd)*2)+(INT(RDAD0_ipd)));

      if (RADDR < 0) then
	RD3_zd := 'X';
	RD2_zd := 'X';
	RD1_zd := 'X';
	RD0_zd := 'X';
	if (TO_X01(RDAD5_ipd) = 'X') and (TO_X01(RDAD5_previous) /= 'X') then
          assert false
	  report ": RDAD5 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD4_ipd) = 'X') and (TO_X01(RDAD4_previous) /= 'X') then
	  assert false
	  report ": RDAD4 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD3_ipd) = 'X') and (TO_X01(RDAD3_previous) /= 'X') then
	  assert false
	  report ": RDAD3 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD2_ipd) = 'X') and (TO_X01(RDAD2_previous) /= 'X') then
	  assert false
	  report ": RDAD2 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD1_ipd) = 'X') and (TO_X01(RDAD1_previous) /= 'X') then
	  assert false
	  report ": RDAD1 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD0_ipd) = 'X') and (TO_X01(RDAD0_previous) /= 'X') then
	  assert false
	  report ": RDAD0 unknown"
	  severity Warning;
	end if;
      else
	RD3_zd := RAM_TMP(RADDR)(3);
	RD2_zd := RAM_TMP(RADDR)(2);
	RD1_zd := RAM_TMP(RADDR)(1);
	RD0_zd := RAM_TMP(RADDR)(0);
      end if;
      
      WCLK_previous := WCLK_ipd;
      WEN_previous := WEN_delayed;
      WEN_delayed := WEN_ipd;
      BLKEN_previous := BLKEN_delayed;
      BLKEN_delayed := BLKEN_ipd;
      WD3_delayed := WD3_ipd;
      WD2_delayed := WD2_ipd;
      WD1_delayed := WD1_ipd;
      WD0_delayed := WD0_ipd;
      WRAD5_previous := WRAD5_delayed;
      WRAD4_previous := WRAD4_delayed;
      WRAD3_previous := WRAD3_delayed;
      WRAD2_previous := WRAD2_delayed;
      WRAD1_previous := WRAD1_delayed;
      WRAD0_previous := WRAD0_delayed;
      WRAD5_delayed := WRAD5_ipd;
      WRAD4_delayed := WRAD4_ipd;
      WRAD3_delayed := WRAD3_ipd;
      WRAD2_delayed := WRAD2_ipd;
      WRAD1_delayed := WRAD1_ipd;
      WRAD0_delayed := WRAD0_ipd;
      RDAD5_previous := RDAD5_ipd;
      RDAD4_previous := RDAD4_ipd;
      RDAD3_previous := RDAD3_ipd;
      RDAD2_previous := RDAD2_ipd;
      RDAD1_previous := RDAD1_ipd;
      RDAD0_previous := RDAD0_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD3,
	GlitchData => RD3_GlitchData,
	OutSignalName => "RD3",
	OutTemp => RD3_zd,
	Paths => (0 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD3), TRUE),
		  1 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
		  2 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
		  3 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
		  4 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  5 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  6 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD3), TRUE),
                  7 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  8 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  9 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  10 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  11 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  12 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD3), TRUE),
                  13 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  14 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  15 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  16 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  17 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  18 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD3), TRUE),
                  19 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  20 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  21 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  22 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  23 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  24 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD3), TRUE),
                  25 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  26 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  27 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  28 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  29 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  30 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD3), TRUE),
                  31 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  32 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  33 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  34 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  35 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD2,
	GlitchData => RD2_GlitchData,
	OutSignalName => "RD2",
	OutTemp => RD2_zd,
	Paths => (0 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD2), TRUE),
		  1 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
		  2 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
		  3 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
		  4 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  5 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  6 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD2), TRUE),
                  7 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  8 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  9 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  10 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  11 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  12 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD2), TRUE),
                  13 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  14 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  15 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  16 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  17 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  18 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD2), TRUE),
                  19 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  20 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  21 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  22 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  23 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  24 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD2), TRUE),
                  25 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  26 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  27 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  28 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  29 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  30 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD2), TRUE),
                  31 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  32 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  33 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  34 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  35 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD1,
	GlitchData => RD1_GlitchData,
	OutSignalName => "RD1",
	OutTemp => RD1_zd,
	Paths => (0 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD1), TRUE),
		  1 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
		  2 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
		  3 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
		  4 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  5 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  6 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD1), TRUE),
                  7 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  8 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  9 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  10 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  11 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  12 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD1), TRUE),
                  13 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  14 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  15 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  16 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  17 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  18 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD1), TRUE),
                  19 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  20 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  21 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  22 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  23 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  24 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD1), TRUE),
                  25 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  26 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  27 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  28 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  29 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  30 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD1), TRUE),
                  31 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  32 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  33 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  34 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  35 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD0,
	GlitchData => RD0_GlitchData,
	OutSignalName => "RD0",
	OutTemp => RD0_zd,
	Paths => (0 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD0), TRUE),
		  1 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
		  2 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
		  3 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
		  4 => (RDAD5_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  5 => (RDAD5_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  6 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD0), TRUE),
                  7 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  8 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  9 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  10 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  11 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  12 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD0), TRUE),
                  13 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  14 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  15 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  16 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  17 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  18 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD0), TRUE),
                  19 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  20 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  21 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  22 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  23 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  24 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD0), TRUE),
                  25 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  26 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  27 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  28 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  29 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  30 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD5_RD0), TRUE),
                  31 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  32 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  33 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  34 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  35 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

  end process VITALBehavior;

end VITAL_ACT;
-----------------------------------------------------------------
--  Proxy Modeling, Inc. 
--
--  Actel RAM4RF VHDL behavioral model
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - Jan/22/96 - Initial Delivery
-- 1.1 - 12/6/96 by DNW - Modified SL_TO_INT.
-- 1.2 - 3/3/97 by DNW - WDx_delayed variables added.
-- 1.3 - 3/6/98 by DNW - Issue "unknown" msg. only if 0/1->X Xtion.
-- 1.4 - 5/27/98 by DNW - Initaialize _ipd signals to X instead of 0.
-- 
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity RAM4RF is
  GENERIC (
        tipd_RDAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD5_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of RAM4RF : entity is TRUE;
  
end RAM4RF;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM4RF is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal WRAD5_ipd : std_ulogic := 'X';
  signal WRAD4_ipd : std_ulogic := 'X';
  signal WRAD3_ipd : std_ulogic := 'X';
  signal WRAD2_ipd : std_ulogic := 'X';
  signal WRAD1_ipd : std_ulogic := 'X';
  signal WRAD0_ipd : std_ulogic := 'X';
  signal WD3_ipd : std_ulogic := 'X';
  signal WD2_ipd : std_ulogic := 'X';
  signal WD1_ipd : std_ulogic := 'X';
  signal WD0_ipd : std_ulogic := 'X';
  signal RDAD5_ipd : std_ulogic := 'X';
  signal RDAD4_ipd : std_ulogic := 'X';
  signal RDAD3_ipd : std_ulogic := 'X';
  signal RDAD2_ipd : std_ulogic := 'X';
  signal RDAD1_ipd : std_ulogic := 'X';
  signal RDAD0_ipd : std_ulogic := 'X';
  signal BLKEN_ipd : std_ulogic := 'X';
  signal WEN_ipd : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal REN_ipd : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  type MEM is array(0 to 63) of std_ulogic_vector(3 downto 0);
   signal RAM_TMP : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (WRAD5_ipd, WRAD5, VitalExtendToFillDelay(tipd_WRAD5));
    VitalWireDelay (WRAD4_ipd, WRAD4, VitalExtendToFillDelay(tipd_WRAD4));
    VitalWireDelay (WRAD3_ipd, WRAD3, VitalExtendToFillDelay(tipd_WRAD3));
    VitalWireDelay (WRAD2_ipd, WRAD2, VitalExtendToFillDelay(tipd_WRAD2));
    VitalWireDelay (WRAD1_ipd, WRAD1, VitalExtendToFillDelay(tipd_WRAD1));
    VitalWireDelay (WRAD0_ipd, WRAD0, VitalExtendToFillDelay(tipd_WRAD0));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (RDAD5_ipd, RDAD5, VitalExtendToFillDelay(tipd_RDAD5));
    VitalWireDelay (RDAD4_ipd, RDAD4, VitalExtendToFillDelay(tipd_RDAD4));
    VitalWireDelay (RDAD3_ipd, RDAD3, VitalExtendToFillDelay(tipd_RDAD3));
    VitalWireDelay (RDAD2_ipd, RDAD2, VitalExtendToFillDelay(tipd_RDAD2));
    VitalWireDelay (RDAD1_ipd, RDAD1, VitalExtendToFillDelay(tipd_RDAD1));
    VitalWireDelay (RDAD0_ipd, RDAD0, VitalExtendToFillDelay(tipd_RDAD0));
    VitalWireDelay (BLKEN_ipd, BLKEN, VitalExtendToFillDelay(tipd_BLKEN));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (REN_ipd, REN, VitalExtendToFillDelay(tipd_REN));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (RDAD5_ipd, RDAD4_ipd, RDAD3_ipd, RDAD2_ipd, 
		RDAD1_ipd, RDAD0_ipd, REN_ipd, RCLK_ipd, 
		WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd, WRAD5_ipd, WRAD4_ipd, 
		WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, WEN_ipd, 
		BLKEN_ipd, BLKENS, WCLK_ipd)

     --  Read Timing Check Results
     variable Tviol_RDAD5_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD5_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD4_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD4_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD3_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD3_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD2_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD2_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD1_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD1_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD0_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD0_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_REN_RCLK_negedge : X01 := '0';
     variable TmDt_REN_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_WD3_WCLK_posedge : X01 := '0';
     variable TmDt_WD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_posedge : X01 := '0';
     variable TmDt_WD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_posedge : X01 := '0';
     variable TmDt_WD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_posedge : X01 := '0';
     variable TmDt_WD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD5_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD4_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD3_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD2_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD1_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD0_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_posedge : X01 := '0';
     variable TmDt_WEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_BLKEN_WCLK_posedge : X01 := '0';
     variable TmDt_BLKEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     --type SL_TO_INT is array(std_ulogic range <>) of integer;
     --constant INT :SL_TO_INT('U' to '-') := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;
  
     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable WEN_delayed : std_ulogic := 'X';
     variable REN_delayed : std_ulogic := 'X';
     variable WEN_previous : std_ulogic := 'X';
     variable REN_previous : std_ulogic := 'X';
     variable BLKEN_delayed : std_ulogic := 'X';
     variable BLKEN_previous : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WRAD5_delayed : std_ulogic := 'X';
     variable WRAD4_delayed : std_ulogic := 'X';
     variable WRAD3_delayed : std_ulogic := 'X';
     variable WRAD2_delayed : std_ulogic := 'X';
     variable WRAD1_delayed : std_ulogic := 'X';
     variable WRAD0_delayed : std_ulogic := 'X';
     variable WRAD5_previous : std_ulogic := 'X';
     variable WRAD4_previous : std_ulogic := 'X';
     variable WRAD3_previous : std_ulogic := 'X';
     variable WRAD2_previous : std_ulogic := 'X';
     variable WRAD1_previous : std_ulogic := 'X';
     variable WRAD0_previous : std_ulogic := 'X';
     variable RDAD5_delayed : std_ulogic := 'X';
     variable RDAD4_delayed : std_ulogic := 'X';
     variable RDAD3_delayed : std_ulogic := 'X';
     variable RDAD2_delayed : std_ulogic := 'X';
     variable RDAD1_delayed : std_ulogic := 'X';
     variable RDAD0_delayed : std_ulogic := 'X';
     variable RDAD5_previous : std_ulogic := 'X';
     variable RDAD4_previous : std_ulogic := 'X';
     variable RDAD3_previous : std_ulogic := 'X';
     variable RDAD2_previous : std_ulogic := 'X';
     variable RDAD1_previous : std_ulogic := 'X';
     variable RDAD0_previous : std_ulogic := 'X';
  
  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RDAD high or low before RCLK falling
      --   Hold  RDAD high or low after RCLK falling

      VitalSetupHoldCheck ( Tviol_RDAD5_RCLK_negedge,
                            TmDt_RDAD5_RCLK_negedge,
                            RDAD5_ipd, "RDAD5",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD5_RCLK_noedge_negedge,
                            tsetup_RDAD5_RCLK_noedge_negedge,
                            thold_RDAD5_RCLK_noedge_negedge,
                            thold_RDAD5_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD4_RCLK_negedge,
                            TmDt_RDAD4_RCLK_negedge,
                            RDAD4_ipd, "RDAD4",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD4_RCLK_noedge_negedge,
                            tsetup_RDAD4_RCLK_noedge_negedge,
                            thold_RDAD4_RCLK_noedge_negedge,
                            thold_RDAD4_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD3_RCLK_negedge,
                            TmDt_RDAD3_RCLK_negedge,
                            RDAD3_ipd, "RDAD3",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD3_RCLK_noedge_negedge,
                            tsetup_RDAD3_RCLK_noedge_negedge,
                            thold_RDAD3_RCLK_noedge_negedge,
                            thold_RDAD3_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD2_RCLK_negedge,
                            TmDt_RDAD2_RCLK_negedge,
                            RDAD2_ipd, "RDAD2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD2_RCLK_noedge_negedge,
                            tsetup_RDAD2_RCLK_noedge_negedge,
                            thold_RDAD2_RCLK_noedge_negedge,
                            thold_RDAD2_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD1_RCLK_negedge,
                            TmDt_RDAD1_RCLK_negedge,
                            RDAD1_ipd, "RDAD1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD1_RCLK_noedge_negedge,
                            tsetup_RDAD1_RCLK_noedge_negedge,
                            thold_RDAD1_RCLK_noedge_negedge,
                            thold_RDAD1_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD0_RCLK_negedge,
                            TmDt_RDAD0_RCLK_negedge,
                            RDAD0_ipd, "RDAD0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD0_RCLK_noedge_negedge,
                            tsetup_RDAD0_RCLK_noedge_negedge,
                            thold_RDAD0_RCLK_noedge_negedge,
                            thold_RDAD0_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup REN high before RCLK falling
      --   Hold  REN high after RCLK falling

      VitalSetupHoldCheck ( Tviol_REN_RCLK_negedge,
                            TmDt_REN_RCLK_negedge,
                            REN_ipd, "REN",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_REN_RCLK_noedge_negedge,
                            tsetup_REN_RCLK_noedge_negedge,
                            thold_REN_RCLK_noedge_negedge,
                            thold_REN_RCLK_noedge_negedge,
                            TimingCheckOn,
                            '\',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup BLKEN high or low before WCLK rising
      --   Hold  BLKEN high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_BLKEN_WCLK_posedge,
                            TmDt_BLKEN_WCLK_posedge,
                            BLKEN_ipd, "BLKEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_BLKEN_WCLK_noedge_posedge,
                            tsetup_BLKEN_WCLK_noedge_posedge,
                            thold_BLKEN_WCLK_noedge_posedge,
                            thold_BLKEN_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WRAD high or low before WCLK rising
      --   Hold  WRAD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WRAD5_WCLK_posedge,
                            TmDt_WRAD5_WCLK_posedge,
                            WRAD5_ipd, "WRAD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD5_WCLK_noedge_posedge,
                            tsetup_WRAD5_WCLK_noedge_posedge,
                            thold_WRAD5_WCLK_noedge_posedge,
                            thold_WRAD5_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD4_WCLK_posedge,
                            TmDt_WRAD4_WCLK_posedge,
                            WRAD4_ipd, "WRAD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD4_WCLK_noedge_posedge,
                            tsetup_WRAD4_WCLK_noedge_posedge,
                            thold_WRAD4_WCLK_noedge_posedge,
                            thold_WRAD4_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD3_WCLK_posedge,
                            TmDt_WRAD3_WCLK_posedge,
                            WRAD3_ipd, "WRAD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD3_WCLK_noedge_posedge,
                            tsetup_WRAD3_WCLK_noedge_posedge,
                            thold_WRAD3_WCLK_noedge_posedge,
                            thold_WRAD3_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD2_WCLK_posedge,
                            TmDt_WRAD2_WCLK_posedge,
                            WRAD2_ipd, "WRAD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD2_WCLK_noedge_posedge,
                            tsetup_WRAD2_WCLK_noedge_posedge,
                            thold_WRAD2_WCLK_noedge_posedge,
                            thold_WRAD2_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD1_WCLK_posedge,
                            TmDt_WRAD1_WCLK_posedge,
                            WRAD1_ipd, "WRAD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD1_WCLK_noedge_posedge,
                            tsetup_WRAD1_WCLK_noedge_posedge,
                            thold_WRAD1_WCLK_noedge_posedge,
                            thold_WRAD1_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD0_WCLK_posedge,
                            TmDt_WRAD0_WCLK_posedge,
                            WRAD0_ipd, "WRAD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD0_WCLK_noedge_posedge,
                            tsetup_WRAD0_WCLK_noedge_posedge,
                            thold_WRAD0_WCLK_noedge_posedge,
                            thold_WRAD0_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WD high or low before WCLK rising
      --   Hold  WD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_posedge,
                            TmDt_WD3_WCLK_posedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_noedge_posedge,
                            tsetup_WD3_WCLK_noedge_posedge,
                            thold_WD3_WCLK_noedge_posedge,
                            thold_WD3_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_posedge,
                            TmDt_WD2_WCLK_posedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_noedge_posedge,
                            tsetup_WD2_WCLK_noedge_posedge,
                            thold_WD2_WCLK_noedge_posedge,
                            thold_WD2_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_posedge,
                            TmDt_WD1_WCLK_posedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_noedge_posedge,
                            tsetup_WD1_WCLK_noedge_posedge,
                            thold_WD1_WCLK_noedge_posedge,
                            thold_WD1_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_posedge,
                            TmDt_WD0_WCLK_posedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_noedge_posedge,
                            tsetup_WD0_WCLK_noedge_posedge,
                            thold_WD0_WCLK_noedge_posedge,
                            thold_WD0_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup WEN high before WCLK rising
      --   Hold  WEN high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_posedge,
                            TmDt_WEN_WCLK_posedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_noedge_posedge,
                            tsetup_WEN_WCLK_noedge_posedge,
                            thold_WEN_WCLK_noedge_posedge,
                            thold_WEN_WCLK_noedge_posedge,
                            (To_X01(BLKEN_ipd)=BLKENS),
                            '/',
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM4RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
    
    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      -- Convert Write Address Signal to Integer
      WADDR := ((INT(WRAD5_delayed)*32)+(INT(WRAD4_delayed)*16)+(INT(WRAD3_delayed)*8)+
		(INT(WRAD2_delayed)*4)+(INT(WRAD1_delayed)*2)+(INT(WRAD0_delayed)));

      if (TO_X01(WCLK_ipd)='X') then
        if (TO_X01(WCLK_previous) /= 'X') then
	  assert false
	  report ": WCLK unknown"
	  severity Warning;
	end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	case TO_X01(WEN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (TO_X01(BLKEN_delayed) = 'X') then
              if (TO_X01(BLKEN_previous) /= 'X') then
	        assert false
	        report ": BLKEN unknown"
	        severity Warning;
	      end if;
	    elsif (TO_X01(BLKEN_delayed) = BLKENS) then
	      if (WADDR < 0) then
		if (TO_X01(WRAD5_delayed) = 'X') and (TO_X01(WRAD5_previous) /= 'X') then
		  assert false
		  report ": WRAD5 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD4_delayed) = 'X') and (TO_X01(WRAD4_previous) /= 'X') then
		  assert false
		  report ": WRAD4 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD3_delayed) = 'X') and (TO_X01(WRAD3_previous) /= 'X') then
		  assert false
		  report ": WRAD3 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD2_delayed) = 'X') and (TO_X01(WRAD2_previous) /= 'X') then
		  assert false
		  report ": WRAD2 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD1_delayed) = 'X') and (TO_X01(WRAD1_previous) /= 'X') then
		  assert false
		  report ": WRAD1 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD0_delayed) = 'X') and (TO_X01(WRAD0_previous) /= 'X') then
		  assert false
		  report ": WRAD0 unknown"
		  severity Warning;
		end if;
	      else 
		RAM_TMP(WADDR) <= WD3_delayed & WD2_delayed & WD1_delayed & WD0_delayed ; 
	      end if;
	    else
	      null;
	    end if;
	  when others =>
            if (TO_X01(WEN_previous) /= 'X') then
	      assert false
	      report ": WEN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      -- Convert Read Address Signal to Integer
      RADDR := ((INT(RDAD5_delayed)*32)+(INT(RDAD4_delayed)*16)+(INT(RDAD3_delayed)*8)+
		(INT(RDAD2_delayed)*4)+(INT(RDAD1_delayed)*2)+(INT(RDAD0_delayed)));

      if (TO_X01(RCLK_ipd) = 'X') then
	RD3_zd := 'X';
	RD2_zd := 'X';
	RD1_zd := 'X';
	RD0_zd := 'X';
	if (TO_X01(RCLK_previous) /= 'X') then
	  assert false
	  report ": RCLK unknown"
	  severity Warning;
	end if;
      elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '0')) then
	case TO_X01(REN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (RADDR < 0) then
	      RD3_zd := 'X';
	      RD2_zd := 'X';
	      RD1_zd := 'X';
	      RD0_zd := 'X';
	      if (TO_X01(RDAD5_delayed) = 'X') and (TO_X01(RDAD5_previous) /= 'X') then
		assert false
		report ": RDAD5 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD4_delayed) = 'X') and (TO_X01(RDAD4_previous) /= 'X') then
		assert false
		report ": RDAD4 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD3_delayed) = 'X') and (TO_X01(RDAD3_previous) /= 'X') then
		assert false
		report ": RDAD3 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD2_delayed) = 'X') and (TO_X01(RDAD2_previous) /= 'X') then
		assert false
		report ": RDAD2 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD1_delayed) = 'X') and (TO_X01(RDAD1_previous) /= 'X') then
		assert false
		report ": RDAD1 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD0_delayed) = 'X') and (TO_X01(RDAD0_previous) /= 'X') then
		assert false
		report ": RDAD0 unknown"
		severity Warning;
	      end if;
	    else
	      RD3_zd := RAM_TMP(RADDR)(3);
	      RD2_zd := RAM_TMP(RADDR)(2);
	      RD1_zd := RAM_TMP(RADDR)(1);
	      RD0_zd := RAM_TMP(RADDR)(0);
	    end if;
	  when others =>
	    RD3_zd := 'X';
	    RD2_zd := 'X';
	    RD1_zd := 'X';
	    RD0_zd := 'X';
            if (TO_X01(REN_previous) /= 'X') then
	      assert false
	      report ": REN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;
      
      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      WEN_previous := WEN_delayed;
      REN_previous := REN_delayed;
      WEN_delayed := WEN_ipd;
      REN_delayed := REN_ipd;
      BLKEN_previous := BLKEN_delayed;
      BLKEN_delayed := BLKEN_ipd;
      WD3_delayed := WD3_ipd;
      WD2_delayed := WD2_ipd;
      WD1_delayed := WD1_ipd;
      WD0_delayed := WD0_ipd;
      WRAD5_previous := WRAD5_delayed;
      WRAD4_previous := WRAD4_delayed;
      WRAD3_previous := WRAD3_delayed;
      WRAD2_previous := WRAD2_delayed;
      WRAD1_previous := WRAD1_delayed;
      WRAD0_previous := WRAD0_delayed;
      WRAD5_delayed := WRAD5_ipd;
      WRAD4_delayed := WRAD4_ipd;
      WRAD3_delayed := WRAD3_ipd;
      WRAD2_delayed := WRAD2_ipd;
      WRAD1_delayed := WRAD1_ipd;
      WRAD0_delayed := WRAD0_ipd;
      RDAD5_previous := RDAD5_delayed;
      RDAD4_previous := RDAD4_delayed;
      RDAD3_previous := RDAD3_delayed;
      RDAD2_previous := RDAD2_delayed;
      RDAD1_previous := RDAD1_delayed;
      RDAD0_previous := RDAD0_delayed;
      RDAD5_delayed := RDAD5_ipd;
      RDAD4_delayed := RDAD4_ipd;
      RDAD3_delayed := RDAD3_ipd;
      RDAD2_delayed := RDAD2_ipd;
      RDAD1_delayed := RDAD1_ipd;
      RDAD0_delayed := RDAD0_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD3,
	GlitchData => RD3_GlitchData,
	OutSignalName => "RD3",
	OutTemp => RD3_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD3), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD2,
	GlitchData => RD2_GlitchData,
	OutSignalName => "RD2",
	OutTemp => RD2_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD2), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD1,
	GlitchData => RD1_GlitchData,
	OutSignalName => "RD1",
	OutTemp => RD1_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD1), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD0,
	GlitchData => RD0_GlitchData,
	OutSignalName => "RD0",
	OutTemp => RD0_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD0), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

  end process VITALBehavior;

end VITAL_ACT;
-----------------------------------------------------------------
--  Proxy Modeling, Inc. 
--
--  Actel RAM4RR VHDL behavioral model
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - Jan/22/96 - Initial Delivery
-- 1.1 - 12/6/96 by DNW - Modified SL_TO_INT.
-- 1.2 - 3/3/97 by DNW - WDx_delayed variables added.
-- 1.3 - 3/6/98 by DNW - Issue "input unknown" msg. only if r/f Xtions.
-- 1.4 - 5/27/98 by DNW - Initaialize _ipd signals to X instead of 0.
-- 
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity RAM4RR is
  GENERIC (
        tipd_RDAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD5    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD5_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD4_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD5_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RDAD5_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD5_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD5  : IN STD_ULOGIC ;
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD5  : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of RAM4RR : entity is TRUE;
  
end RAM4RR;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM4RR is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal WRAD5_ipd : std_ulogic := 'X';
  signal WRAD4_ipd : std_ulogic := 'X';
  signal WRAD3_ipd : std_ulogic := 'X';
  signal WRAD2_ipd : std_ulogic := 'X';
  signal WRAD1_ipd : std_ulogic := 'X';
  signal WRAD0_ipd : std_ulogic := 'X';
  signal WD3_ipd : std_ulogic := 'X';
  signal WD2_ipd : std_ulogic := 'X';
  signal WD1_ipd : std_ulogic := 'X';
  signal WD0_ipd : std_ulogic := 'X';
  signal RDAD5_ipd : std_ulogic := 'X';
  signal RDAD4_ipd : std_ulogic := 'X';
  signal RDAD3_ipd : std_ulogic := 'X';
  signal RDAD2_ipd : std_ulogic := 'X';
  signal RDAD1_ipd : std_ulogic := 'X';
  signal RDAD0_ipd : std_ulogic := 'X';
  signal BLKEN_ipd : std_ulogic := 'X';
  signal WEN_ipd : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal REN_ipd : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  type MEM is array(0 to 63) of std_ulogic_vector(3 downto 0);
   signal RAM_TMP : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (WRAD5_ipd, WRAD5, VitalExtendToFillDelay(tipd_WRAD5));
    VitalWireDelay (WRAD4_ipd, WRAD4, VitalExtendToFillDelay(tipd_WRAD4));
    VitalWireDelay (WRAD3_ipd, WRAD3, VitalExtendToFillDelay(tipd_WRAD3));
    VitalWireDelay (WRAD2_ipd, WRAD2, VitalExtendToFillDelay(tipd_WRAD2));
    VitalWireDelay (WRAD1_ipd, WRAD1, VitalExtendToFillDelay(tipd_WRAD1));
    VitalWireDelay (WRAD0_ipd, WRAD0, VitalExtendToFillDelay(tipd_WRAD0));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (RDAD5_ipd, RDAD5, VitalExtendToFillDelay(tipd_RDAD5));
    VitalWireDelay (RDAD4_ipd, RDAD4, VitalExtendToFillDelay(tipd_RDAD4));
    VitalWireDelay (RDAD3_ipd, RDAD3, VitalExtendToFillDelay(tipd_RDAD3));
    VitalWireDelay (RDAD2_ipd, RDAD2, VitalExtendToFillDelay(tipd_RDAD2));
    VitalWireDelay (RDAD1_ipd, RDAD1, VitalExtendToFillDelay(tipd_RDAD1));
    VitalWireDelay (RDAD0_ipd, RDAD0, VitalExtendToFillDelay(tipd_RDAD0));
    VitalWireDelay (BLKEN_ipd, BLKEN, VitalExtendToFillDelay(tipd_BLKEN));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (REN_ipd, REN, VitalExtendToFillDelay(tipd_REN));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (RDAD5_ipd, RDAD4_ipd, RDAD3_ipd, RDAD2_ipd, 
		RDAD1_ipd, RDAD0_ipd, REN_ipd, RCLK_ipd, 
		WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd, WRAD5_ipd, WRAD4_ipd, 
		WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, WEN_ipd, 
		BLKEN_ipd, BLKENS, WCLK_ipd)

     --  Read Timing Check Results
     variable Tviol_RDAD5_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD5_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD4_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD4_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD3_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD2_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD1_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD0_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_REN_RCLK_posedge : X01 := '0';
     variable TmDt_REN_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_WD3_WCLK_posedge : X01 := '0';
     variable TmDt_WD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_posedge : X01 := '0';
     variable TmDt_WD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_posedge : X01 := '0';
     variable TmDt_WD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_posedge : X01 := '0';
     variable TmDt_WD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD5_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD4_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD3_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD2_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD1_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD0_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_posedge : X01 := '0';
     variable TmDt_WEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_BLKEN_WCLK_posedge : X01 := '0';
     variable TmDt_BLKEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     --type SL_TO_INT is array(std_ulogic range <>) of integer;
     --constant INT :SL_TO_INT('U' to '-') := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;

     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable WEN_delayed : std_ulogic := 'X';
     variable REN_delayed : std_ulogic := 'X';
     variable WEN_previous : std_ulogic := 'X';
     variable REN_previous : std_ulogic := 'X';
     variable BLKEN_delayed : std_ulogic := 'X';
     variable BLKEN_previous : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WRAD5_delayed : std_ulogic := 'X';
     variable WRAD4_delayed : std_ulogic := 'X';
     variable WRAD3_delayed : std_ulogic := 'X';
     variable WRAD2_delayed : std_ulogic := 'X';
     variable WRAD1_delayed : std_ulogic := 'X';
     variable WRAD0_delayed : std_ulogic := 'X';
     variable WRAD5_previous : std_ulogic := 'X';
     variable WRAD4_previous : std_ulogic := 'X';
     variable WRAD3_previous : std_ulogic := 'X';
     variable WRAD2_previous : std_ulogic := 'X';
     variable WRAD1_previous : std_ulogic := 'X';
     variable WRAD0_previous : std_ulogic := 'X';
     variable RDAD5_delayed : std_ulogic := 'X';
     variable RDAD4_delayed : std_ulogic := 'X';
     variable RDAD3_delayed : std_ulogic := 'X';
     variable RDAD2_delayed : std_ulogic := 'X';
     variable RDAD1_delayed : std_ulogic := 'X';
     variable RDAD0_delayed : std_ulogic := 'X';
     variable RDAD5_previous : std_ulogic := 'X';
     variable RDAD4_previous : std_ulogic := 'X';
     variable RDAD3_previous : std_ulogic := 'X';
     variable RDAD2_previous : std_ulogic := 'X';
     variable RDAD1_previous : std_ulogic := 'X';
     variable RDAD0_previous : std_ulogic := 'X';
  
  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RDAD high or low before RCLK rising
      --   Hold  RDAD high or low after RCLK rising

      VitalSetupHoldCheck ( Tviol_RDAD5_RCLK_posedge,
                            TmDt_RDAD5_RCLK_posedge,
                            RDAD5_ipd, "RDAD5",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD5_RCLK_noedge_posedge,
                            tsetup_RDAD5_RCLK_noedge_posedge,
                            thold_RDAD5_RCLK_noedge_posedge,
                            thold_RDAD5_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD4_RCLK_posedge,
                            TmDt_RDAD4_RCLK_posedge,
                            RDAD4_ipd, "RDAD4",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD4_RCLK_noedge_posedge,
                            tsetup_RDAD4_RCLK_noedge_posedge,
                            thold_RDAD4_RCLK_noedge_posedge,
                            thold_RDAD4_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD3_RCLK_posedge,
                            TmDt_RDAD3_RCLK_posedge,
                            RDAD3_ipd, "RDAD3",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD3_RCLK_noedge_posedge,
                            tsetup_RDAD3_RCLK_noedge_posedge,
                            thold_RDAD3_RCLK_noedge_posedge,
                            thold_RDAD3_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD2_RCLK_posedge,
                            TmDt_RDAD2_RCLK_posedge,
                            RDAD2_ipd, "RDAD2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD2_RCLK_noedge_posedge,
                            tsetup_RDAD2_RCLK_noedge_posedge,
                            thold_RDAD2_RCLK_noedge_posedge,
                            thold_RDAD2_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD1_RCLK_posedge,
                            TmDt_RDAD1_RCLK_posedge,
                            RDAD1_ipd, "RDAD1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD1_RCLK_noedge_posedge,
                            tsetup_RDAD1_RCLK_noedge_posedge,
                            thold_RDAD1_RCLK_noedge_posedge,
                            thold_RDAD1_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD0_RCLK_posedge,
                            TmDt_RDAD0_RCLK_posedge,
                            RDAD0_ipd, "RDAD0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD0_RCLK_noedge_posedge,
                            tsetup_RDAD0_RCLK_noedge_posedge,
                            thold_RDAD0_RCLK_noedge_posedge,
                            thold_RDAD0_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup REN high before RCLK rising
      --   Hold  REN high after RCLK rising

      VitalSetupHoldCheck ( Tviol_REN_RCLK_posedge,
                            TmDt_REN_RCLK_posedge,
                            REN_ipd, "REN",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_REN_RCLK_noedge_posedge,
                            tsetup_REN_RCLK_noedge_posedge,
                            thold_REN_RCLK_noedge_posedge,
                            thold_REN_RCLK_noedge_posedge,
                            TimingCheckOn,
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup BLKEN high or low before WCLK rising
      --   Hold  BLKEN high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_BLKEN_WCLK_posedge,
                            TmDt_BLKEN_WCLK_posedge,
                            BLKEN_ipd, "BLKEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_BLKEN_WCLK_noedge_posedge,
                            tsetup_BLKEN_WCLK_noedge_posedge,
                            thold_BLKEN_WCLK_noedge_posedge,
                            thold_BLKEN_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WRAD high or low before WCLK rising
      --   Hold  WRAD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WRAD5_WCLK_posedge,
                            TmDt_WRAD5_WCLK_posedge,
                            WRAD5_ipd, "WRAD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD5_WCLK_noedge_posedge,
                            tsetup_WRAD5_WCLK_noedge_posedge,
                            thold_WRAD5_WCLK_noedge_posedge,
                            thold_WRAD5_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD4_WCLK_posedge,
                            TmDt_WRAD4_WCLK_posedge,
                            WRAD4_ipd, "WRAD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD4_WCLK_noedge_posedge,
                            tsetup_WRAD4_WCLK_noedge_posedge,
                            thold_WRAD4_WCLK_noedge_posedge,
                            thold_WRAD4_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD3_WCLK_posedge,
                            TmDt_WRAD3_WCLK_posedge,
                            WRAD3_ipd, "WRAD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD3_WCLK_noedge_posedge,
                            tsetup_WRAD3_WCLK_noedge_posedge,
                            thold_WRAD3_WCLK_noedge_posedge,
                            thold_WRAD3_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD2_WCLK_posedge,
                            TmDt_WRAD2_WCLK_posedge,
                            WRAD2_ipd, "WRAD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD2_WCLK_noedge_posedge,
                            tsetup_WRAD2_WCLK_noedge_posedge,
                            thold_WRAD2_WCLK_noedge_posedge,
                            thold_WRAD2_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD1_WCLK_posedge,
                            TmDt_WRAD1_WCLK_posedge,
                            WRAD1_ipd, "WRAD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD1_WCLK_noedge_posedge,
                            tsetup_WRAD1_WCLK_noedge_posedge,
                            thold_WRAD1_WCLK_noedge_posedge,
                            thold_WRAD1_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD0_WCLK_posedge,
                            TmDt_WRAD0_WCLK_posedge,
                            WRAD0_ipd, "WRAD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD0_WCLK_noedge_posedge,
                            tsetup_WRAD0_WCLK_noedge_posedge,
                            thold_WRAD0_WCLK_noedge_posedge,
                            thold_WRAD0_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WD high or low before WCLK rising
      --   Hold  WD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_posedge,
                            TmDt_WD3_WCLK_posedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_noedge_posedge,
                            tsetup_WD3_WCLK_noedge_posedge,
                            thold_WD3_WCLK_noedge_posedge,
                            thold_WD3_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_posedge,
                            TmDt_WD2_WCLK_posedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_noedge_posedge,
                            tsetup_WD2_WCLK_noedge_posedge,
                            thold_WD2_WCLK_noedge_posedge,
                            thold_WD2_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_posedge,
                            TmDt_WD1_WCLK_posedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_noedge_posedge,
                            tsetup_WD1_WCLK_noedge_posedge,
                            thold_WD1_WCLK_noedge_posedge,
                            thold_WD1_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_posedge,
                            TmDt_WD0_WCLK_posedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_noedge_posedge,
                            tsetup_WD0_WCLK_noedge_posedge,
                            thold_WD0_WCLK_noedge_posedge,
                            thold_WD0_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup WEN high before WCLK rising
      --   Hold  WEN high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_posedge,
                            TmDt_WEN_WCLK_posedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_noedge_posedge,
                            tsetup_WEN_WCLK_noedge_posedge,
                            thold_WEN_WCLK_noedge_posedge,
                            thold_WEN_WCLK_noedge_posedge,
                            (To_X01(BLKEN_ipd)=BLKENS),
                            '/',
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM4RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
    
    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      -- Convert Write Address Signal to Integer
      WADDR := ((INT(WRAD5_delayed)*32)+(INT(WRAD4_delayed)*16)+(INT(WRAD3_delayed)*8)+
		(INT(WRAD2_delayed)*4)+(INT(WRAD1_delayed)*2)+(INT(WRAD0_delayed)));

      if (TO_X01(WCLK_ipd)='X') then
        if (TO_X01(WCLK_previous) /= 'X') then
	  assert false
	  report ": WCLK unknown"
	  severity Warning;
	end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	case TO_X01(WEN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (TO_X01(BLKEN_delayed) = 'X') then
              if (TO_X01(BLKEN_previous) /= 'X') then
	        assert false
	        report ": BLKEN unknown"
	        severity Warning;
	      end if;
	    elsif (TO_X01(BLKEN_delayed) = BLKENS) then
	      if (WADDR < 0) then
		if (TO_X01(WRAD5_delayed) = 'X') and (TO_X01(WRAD5_previous) /= 'X') then
		  assert false
		  report ": WRAD5 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD4_delayed) = 'X') and (TO_X01(WRAD4_previous) /= 'X') then
		  assert false
		  report ": WRAD4 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD3_delayed) = 'X') and (TO_X01(WRAD3_previous) /= 'X') then
		  assert false
		  report ": WRAD3 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD2_delayed) = 'X') and (TO_X01(WRAD2_previous) /= 'X') then
		  assert false
		  report ": WRAD2 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD1_delayed) = 'X') and (TO_X01(WRAD1_previous) /= 'X') then
		  assert false
		  report ": WRAD1 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD0_delayed) = 'X') and (TO_X01(WRAD0_previous) /= 'X') then
		  assert false
		  report ": WRAD0 unknown"
		  severity Warning;
		end if;
	      else 
		RAM_TMP(WADDR) <= WD3_delayed & WD2_delayed & WD1_delayed & WD0_delayed ; 
	      end if;
	    else
	      null;
	    end if;
	  when others =>
            if (TO_X01(WEN_previous) /= 'X') then
	      assert false
	      report ": WEN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      -- Convert Read Address Signal to Integer
      RADDR := ((INT(RDAD5_delayed)*32)+(INT(RDAD4_delayed)*16)+(INT(RDAD3_delayed)*8)+
		(INT(RDAD2_delayed)*4)+(INT(RDAD1_delayed)*2)+(INT(RDAD0_delayed)));

      if (TO_X01(RCLK_ipd) = 'X') then
	RD3_zd := 'X';
	RD2_zd := 'X';
	RD1_zd := 'X';
	RD0_zd := 'X';
	if (TO_X01(RCLK_previous) /= 'X') then
	  assert false
	  report ": RCLK unknown"
	  severity Warning;
	end if;
      elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1')) then
	case TO_X01(REN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (RADDR < 0) then
	      RD3_zd := 'X';
	      RD2_zd := 'X';
	      RD1_zd := 'X';
	      RD0_zd := 'X';
	      if (TO_X01(RDAD5_delayed) = 'X') and (TO_X01(RDAD5_previous) /= 'X') then
		assert false
		report ": RDAD5 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD4_delayed) = 'X') and (TO_X01(RDAD4_previous) /= 'X') then
		assert false
		report ": RDAD4 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD3_delayed) = 'X') and (TO_X01(RDAD3_previous) /= 'X') then
		assert false
		report ": RDAD3 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD2_delayed) = 'X') and (TO_X01(RDAD2_previous) /= 'X') then
		assert false
		report ": RDAD2 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD1_delayed) = 'X') and (TO_X01(RDAD1_previous) /= 'X') then
		assert false
		report ": RDAD1 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD0_delayed) = 'X') and (TO_X01(RDAD0_previous) /= 'X') then
		assert false
		report ": RDAD0 unknown"
		severity Warning;
	      end if;
	    else
	      RD3_zd := RAM_TMP(RADDR)(3);
	      RD2_zd := RAM_TMP(RADDR)(2);
	      RD1_zd := RAM_TMP(RADDR)(1);
	      RD0_zd := RAM_TMP(RADDR)(0);
	    end if;
	  when others =>
	    RD3_zd := 'X';
	    RD2_zd := 'X';
	    RD1_zd := 'X';
	    RD0_zd := 'X';
            if (TO_X01(REN_previous) /= 'X') then
	      assert false
	      report ": REN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;
      
      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      WEN_previous := WEN_delayed;
      REN_previous := REN_delayed;
      WEN_delayed := WEN_ipd;
      REN_delayed := REN_ipd;
      BLKEN_previous := BLKEN_delayed;
      BLKEN_delayed := BLKEN_ipd;
      WD3_delayed := WD3_ipd;
      WD2_delayed := WD2_ipd;
      WD1_delayed := WD1_ipd;
      WD0_delayed := WD0_ipd;
      WRAD5_previous := WRAD5_delayed;
      WRAD4_previous := WRAD4_delayed;
      WRAD3_previous := WRAD3_delayed;
      WRAD2_previous := WRAD2_delayed;
      WRAD1_previous := WRAD1_delayed;
      WRAD0_previous := WRAD0_delayed;
      WRAD5_delayed := WRAD5_ipd;
      WRAD4_delayed := WRAD4_ipd;
      WRAD3_delayed := WRAD3_ipd;
      WRAD2_delayed := WRAD2_ipd;
      WRAD1_delayed := WRAD1_ipd;
      WRAD0_delayed := WRAD0_ipd;
      RDAD5_previous := RDAD5_delayed;
      RDAD4_previous := RDAD4_delayed;
      RDAD3_previous := RDAD3_delayed;
      RDAD2_previous := RDAD2_delayed;
      RDAD1_previous := RDAD1_delayed;
      RDAD0_previous := RDAD0_delayed;
      RDAD5_delayed := RDAD5_ipd;
      RDAD4_delayed := RDAD4_ipd;
      RDAD3_delayed := RDAD3_ipd;
      RDAD2_delayed := RDAD2_ipd;
      RDAD1_delayed := RDAD1_ipd;
      RDAD0_delayed := RDAD0_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD3,
	GlitchData => RD3_GlitchData,
	OutSignalName => "RD3",
	OutTemp => RD3_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD3), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD2,
	GlitchData => RD2_GlitchData,
	OutSignalName => "RD2",
	OutTemp => RD2_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD2), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD1,
	GlitchData => RD1_GlitchData,
	OutSignalName => "RD1",
	OutTemp => RD1_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD1), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD0,
	GlitchData => RD0_GlitchData,
	OutSignalName => "RD0",
	OutTemp => RD0_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD0), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

  end process VITALBehavior;

end VITAL_ACT;
-----------------------------------------------------------------
--  Proxy Modeling, Inc. 
--
--  Actel RAM8FA VHDL behavioral model
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - Jan/22/96 - Initial Delivery
-- 1.1 - 12/6/96 by DNW - Modified SL_TO_INT.
-- 1.2 - 3/3/97 by DNW - WDx_delayed variables added.
-- 1.3 - 3/6/98 by DNW - Issue "unknown" msg. only if 0/1->X Xtion.
-- 1.4 - 5/27/98 by DNW - Initaialize _ipd signals to X instead of 0.
-- 
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity RAM8FA is
  GENERIC (
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD7      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD6      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD5      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD4      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RDAD4_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_WRAD4_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC;
        RD6    : OUT STD_ULOGIC;
        RD5    : OUT STD_ULOGIC;
        RD4    : OUT STD_ULOGIC;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of RAM8FA : entity is TRUE;
  
end RAM8FA;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM8FA is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal WRAD4_ipd : std_ulogic := 'X';
  signal WRAD3_ipd : std_ulogic := 'X';
  signal WRAD2_ipd : std_ulogic := 'X';
  signal WRAD1_ipd : std_ulogic := 'X';
  signal WRAD0_ipd : std_ulogic := 'X';
  signal WD7_ipd : std_ulogic := 'X';
  signal WD6_ipd : std_ulogic := 'X';
  signal WD5_ipd : std_ulogic := 'X';
  signal WD4_ipd : std_ulogic := 'X';
  signal WD3_ipd : std_ulogic := 'X';
  signal WD2_ipd : std_ulogic := 'X';
  signal WD1_ipd : std_ulogic := 'X';
  signal WD0_ipd : std_ulogic := 'X';
  signal RDAD4_ipd : std_ulogic := 'X';
  signal RDAD3_ipd : std_ulogic := 'X';
  signal RDAD2_ipd : std_ulogic := 'X';
  signal RDAD1_ipd : std_ulogic := 'X';
  signal RDAD0_ipd : std_ulogic := 'X';
  signal BLKEN_ipd : std_ulogic := 'X';
  signal WEN_ipd : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  type MEM is array(0 to 31) of std_ulogic_vector(7 downto 0);
   signal RAM_TMP : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (WRAD4_ipd, WRAD4, VitalExtendToFillDelay(tipd_WRAD4));
    VitalWireDelay (WRAD3_ipd, WRAD3, VitalExtendToFillDelay(tipd_WRAD3));
    VitalWireDelay (WRAD2_ipd, WRAD2, VitalExtendToFillDelay(tipd_WRAD2));
    VitalWireDelay (WRAD1_ipd, WRAD1, VitalExtendToFillDelay(tipd_WRAD1));
    VitalWireDelay (WRAD0_ipd, WRAD0, VitalExtendToFillDelay(tipd_WRAD0));
    VitalWireDelay (WD7_ipd, WD7, VitalExtendToFillDelay(tipd_WD7));
    VitalWireDelay (WD6_ipd, WD6, VitalExtendToFillDelay(tipd_WD6));
    VitalWireDelay (WD5_ipd, WD5, VitalExtendToFillDelay(tipd_WD5));
    VitalWireDelay (WD4_ipd, WD4, VitalExtendToFillDelay(tipd_WD4));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (RDAD4_ipd, RDAD4, VitalExtendToFillDelay(tipd_RDAD4));
    VitalWireDelay (RDAD3_ipd, RDAD3, VitalExtendToFillDelay(tipd_RDAD3));
    VitalWireDelay (RDAD2_ipd, RDAD2, VitalExtendToFillDelay(tipd_RDAD2));
    VitalWireDelay (RDAD1_ipd, RDAD1, VitalExtendToFillDelay(tipd_RDAD1));
    VitalWireDelay (RDAD0_ipd, RDAD0, VitalExtendToFillDelay(tipd_RDAD0));
    VitalWireDelay (BLKEN_ipd, BLKEN, VitalExtendToFillDelay(tipd_BLKEN));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (RDAD4_ipd, RDAD3_ipd, RDAD2_ipd, RDAD1_ipd, 
		RDAD0_ipd, WD7_ipd, WD6_ipd, WD5_ipd, 
		WD4_ipd, WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd, WRAD4_ipd, 
		WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, WEN_ipd, 
		BLKEN_ipd, BLKENS, WCLK_ipd, RAM_TMP)

     --  Write Timing Check Results
     variable Tviol_WD7_WCLK_negedge : X01 := '0';
     variable TmDt_WD7_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD6_WCLK_negedge : X01 := '0';
     variable TmDt_WD6_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD5_WCLK_negedge : X01 := '0';
     variable TmDt_WD5_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD4_WCLK_negedge : X01 := '0';
     variable TmDt_WD4_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD3_WCLK_negedge : X01 := '0';
     variable TmDt_WD3_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_negedge : X01 := '0';
     variable TmDt_WD2_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_negedge : X01 := '0';
     variable TmDt_WD1_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_negedge : X01 := '0';
     variable TmDt_WD0_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD4_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD4_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD3_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD3_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD2_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD2_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD1_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD1_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD0_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD0_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_negedge : X01 := '0';
     variable TmDt_WEN_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_BLKEN_WCLK_negedge : X01 := '0';
     variable TmDt_BLKEN_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     --type SL_TO_INT is array(std_ulogic range <>) of integer;
     --constant INT :SL_TO_INT('U' to '-') := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     variable RD7_zd : std_ulogic;
     variable RD6_zd : std_ulogic;
     variable RD5_zd : std_ulogic;
     variable RD4_zd : std_ulogic;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD7_GlitchData : VitalGlitchDataType;
     variable RD6_GlitchData : VitalGlitchDataType;
     variable RD5_GlitchData : VitalGlitchDataType;
     variable RD4_GlitchData : VitalGlitchDataType;
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;
  
     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable WEN_delayed : std_ulogic := 'X';
     variable WEN_previous : std_ulogic := 'X';
     variable BLKEN_delayed : std_ulogic := 'X';
     variable BLKEN_previous : std_ulogic := 'X';
     variable WD7_delayed : std_ulogic := 'X';
     variable WD6_delayed : std_ulogic := 'X';
     variable WD5_delayed : std_ulogic := 'X';
     variable WD4_delayed : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WRAD4_delayed : std_ulogic := 'X';
     variable WRAD3_delayed : std_ulogic := 'X';
     variable WRAD2_delayed : std_ulogic := 'X';
     variable WRAD1_delayed : std_ulogic := 'X';
     variable WRAD0_delayed : std_ulogic := 'X';
     variable WRAD4_previous : std_ulogic := 'X';
     variable WRAD3_previous : std_ulogic := 'X';
     variable WRAD2_previous : std_ulogic := 'X';
     variable WRAD1_previous : std_ulogic := 'X';
     variable WRAD0_previous : std_ulogic := 'X';
     variable RDAD4_previous : std_ulogic := 'X';
     variable RDAD3_previous : std_ulogic := 'X';
     variable RDAD2_previous : std_ulogic := 'X';
     variable RDAD1_previous : std_ulogic := 'X';
     variable RDAD0_previous : std_ulogic := 'X';
  
  begin  --  process VITALBehavior 

    if (TimingCheckOn) then

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup BLKEN high or low before WCLK falling
      --   Hold  BLKEN high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_BLKEN_WCLK_negedge,
                            TmDt_BLKEN_WCLK_negedge,
                            BLKEN_ipd, "BLKEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_BLKEN_WCLK_noedge_negedge,
                            tsetup_BLKEN_WCLK_noedge_negedge,
                            thold_BLKEN_WCLK_noedge_negedge,
                            thold_BLKEN_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WRAD high or low before WCLK falling
      --   Hold  WRAD high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_WRAD4_WCLK_negedge,
                            TmDt_WRAD4_WCLK_negedge,
                            WRAD4_ipd, "WRAD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD4_WCLK_noedge_negedge,
                            tsetup_WRAD4_WCLK_noedge_negedge,
                            thold_WRAD4_WCLK_noedge_negedge,
                            thold_WRAD4_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD3_WCLK_negedge,
                            TmDt_WRAD3_WCLK_negedge,
                            WRAD3_ipd, "WRAD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD3_WCLK_noedge_negedge,
                            tsetup_WRAD3_WCLK_noedge_negedge,
                            thold_WRAD3_WCLK_noedge_negedge,
                            thold_WRAD3_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD2_WCLK_negedge,
                            TmDt_WRAD2_WCLK_negedge,
                            WRAD2_ipd, "WRAD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD2_WCLK_noedge_negedge,
                            tsetup_WRAD2_WCLK_noedge_negedge,
                            thold_WRAD2_WCLK_noedge_negedge,
                            thold_WRAD2_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD1_WCLK_negedge,
                            TmDt_WRAD1_WCLK_negedge,
                            WRAD1_ipd, "WRAD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD1_WCLK_noedge_negedge,
                            tsetup_WRAD1_WCLK_noedge_negedge,
                            thold_WRAD1_WCLK_noedge_negedge,
                            thold_WRAD1_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD0_WCLK_negedge,
                            TmDt_WRAD0_WCLK_negedge,
                            WRAD0_ipd, "WRAD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD0_WCLK_noedge_negedge,
                            tsetup_WRAD0_WCLK_noedge_negedge,
                            thold_WRAD0_WCLK_noedge_negedge,
                            thold_WRAD0_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WD high or low before WCLK falling
      --   Hold  WD high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_WD7_WCLK_negedge,
                            TmDt_WD7_WCLK_negedge,
                            WD7_ipd, "WD7",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD7_WCLK_noedge_negedge,
                            tsetup_WD7_WCLK_noedge_negedge,
                            thold_WD7_WCLK_noedge_negedge,
                            thold_WD7_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD6_WCLK_negedge,
                            TmDt_WD6_WCLK_negedge,
                            WD6_ipd, "WD6",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD6_WCLK_noedge_negedge,
                            tsetup_WD6_WCLK_noedge_negedge,
                            thold_WD6_WCLK_noedge_negedge,
                            thold_WD6_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD5_WCLK_negedge,
                            TmDt_WD5_WCLK_negedge,
                            WD5_ipd, "WD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD5_WCLK_noedge_negedge,
                            tsetup_WD5_WCLK_noedge_negedge,
                            thold_WD5_WCLK_noedge_negedge,
                            thold_WD5_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD4_WCLK_negedge,
                            TmDt_WD4_WCLK_negedge,
                            WD4_ipd, "WD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD4_WCLK_noedge_negedge,
                            tsetup_WD4_WCLK_noedge_negedge,
                            thold_WD4_WCLK_noedge_negedge,
                            thold_WD4_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_negedge,
                            TmDt_WD3_WCLK_negedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_noedge_negedge,
                            tsetup_WD3_WCLK_noedge_negedge,
                            thold_WD3_WCLK_noedge_negedge,
                            thold_WD3_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_negedge,
                            TmDt_WD2_WCLK_negedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_noedge_negedge,
                            tsetup_WD2_WCLK_noedge_negedge,
                            thold_WD2_WCLK_noedge_negedge,
                            thold_WD2_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_negedge,
                            TmDt_WD1_WCLK_negedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_noedge_negedge,
                            tsetup_WD1_WCLK_noedge_negedge,
                            thold_WD1_WCLK_noedge_negedge,
                            thold_WD1_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_negedge,
                            TmDt_WD0_WCLK_negedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_noedge_negedge,
                            tsetup_WD0_WCLK_noedge_negedge,
                            thold_WD0_WCLK_noedge_negedge,
                            thold_WD0_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup WEN high before WCLK falling
      --   Hold  WEN high after WCLK falling

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_negedge,
                            TmDt_WEN_WCLK_negedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_noedge_negedge,
                            tsetup_WEN_WCLK_noedge_negedge,
                            thold_WEN_WCLK_noedge_negedge,
                            thold_WEN_WCLK_noedge_negedge,
                            (To_X01(BLKEN_ipd)=BLKENS),
                            '\',
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM8FA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
    
    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      -- Convert Write Address Signal to Integer
      WADDR := ((INT(WRAD4_delayed)*16)+(INT(WRAD3_delayed)*8)+(INT(WRAD2_delayed)*4)
		+(INT(WRAD1_delayed)*2)+(INT(WRAD0_delayed)));

      if (TO_X01(WCLK_ipd)='X') then
        if (TO_X01(WCLK_previous) /= 'X') then
	  assert false
	  report ": WCLK unknown"
	  severity Warning;
	end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='0')) then
	case TO_X01(WEN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (TO_X01(BLKEN_delayed) = 'X') then
              if (TO_X01(BLKEN_previous) /= 'X') then
	        assert false
	        report ": BLKEN unknown"
	        severity Warning;
	      end if;
	    elsif (TO_X01(BLKEN_delayed) = BLKENS) then
	      if (WADDR < 0) then
		if (TO_X01(WRAD4_delayed) = 'X') and (TO_X01(WRAD4_previous) /= 'X') then
		  assert false
		  report ": WRAD4 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD3_delayed) = 'X') and (TO_X01(WRAD3_previous) /= 'X') then
		  assert false
		  report ": WRAD3 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD2_delayed) = 'X') and (TO_X01(WRAD2_previous) /= 'X') then
		  assert false
		  report ": WRAD2 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD1_delayed) = 'X') and (TO_X01(WRAD1_previous) /= 'X') then
		  assert false
		  report ": WRAD1 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD0_delayed) = 'X') and (TO_X01(WRAD0_previous) /= 'X') then
		  assert false
		  report ": WRAD0 unknown"
		  severity Warning;
		end if;
	      else 
		RAM_TMP(WADDR) <= WD7_delayed & WD6_delayed & WD5_delayed & 
                                  WD4_delayed & WD3_delayed & WD2_delayed &
                                  WD1_delayed & WD0_delayed ; 
	      end if;
	    else
	      null;
	    end if;
	  when others =>
            if (TO_X01(WEN_previous) /= 'X') then
	      assert false
	      report ": WEN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      -- Convert Read Address Signal to Integer
      RADDR := ((INT(RDAD4_ipd)*16)+(INT(RDAD3_ipd)*8)+
		(INT(RDAD2_ipd)*4)+(INT(RDAD1_ipd)*2)+(INT(RDAD0_ipd)));

      if (RADDR < 0) then
	RD7_zd := 'X';
	RD6_zd := 'X';
	RD5_zd := 'X';
	RD4_zd := 'X';
	RD3_zd := 'X';
	RD2_zd := 'X';
	RD1_zd := 'X';
	RD0_zd := 'X';
	if (TO_X01(RDAD4_ipd) = 'X') and (TO_X01(RDAD4_previous) /= 'X') then
	  assert false
	  report ": RDAD4 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD3_ipd) = 'X') and (TO_X01(RDAD3_previous) /= 'X') then
	  assert false
	  report ": RDAD3 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD2_ipd) = 'X') and (TO_X01(RDAD2_previous) /= 'X') then
	  assert false
	  report ": RDAD2 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD1_ipd) = 'X') and (TO_X01(RDAD1_previous) /= 'X') then
	  assert false
	  report ": RDAD1 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD0_ipd) = 'X') and (TO_X01(RDAD0_previous) /= 'X') then
	  assert false
	  report ": RDAD0 unknown"
	  severity Warning;
	end if;
      else
	RD7_zd := RAM_TMP(RADDR)(7);
	RD6_zd := RAM_TMP(RADDR)(6);
	RD5_zd := RAM_TMP(RADDR)(5);
	RD4_zd := RAM_TMP(RADDR)(4);
	RD3_zd := RAM_TMP(RADDR)(3);
	RD2_zd := RAM_TMP(RADDR)(2);
	RD1_zd := RAM_TMP(RADDR)(1);
	RD0_zd := RAM_TMP(RADDR)(0);
      end if;
      
      WCLK_previous := WCLK_ipd;
      WEN_previous := WEN_delayed;
      WEN_delayed := WEN_ipd;
      BLKEN_previous := BLKEN_delayed;
      BLKEN_delayed := BLKEN_ipd;
      WD7_delayed := WD7_ipd;
      WD6_delayed := WD6_ipd;
      WD5_delayed := WD5_ipd;
      WD4_delayed := WD4_ipd;
      WD3_delayed := WD3_ipd;
      WD2_delayed := WD2_ipd;
      WD1_delayed := WD1_ipd;
      WD0_delayed := WD0_ipd;
      WRAD4_previous := WRAD4_delayed;
      WRAD3_previous := WRAD3_delayed;
      WRAD2_previous := WRAD2_delayed;
      WRAD1_previous := WRAD1_delayed;
      WRAD0_previous := WRAD0_delayed;
      WRAD4_delayed := WRAD4_ipd;
      WRAD3_delayed := WRAD3_ipd;
      WRAD2_delayed := WRAD2_ipd;
      WRAD1_delayed := WRAD1_ipd;
      WRAD0_delayed := WRAD0_ipd;
      RDAD4_previous := RDAD4_ipd;
      RDAD3_previous := RDAD3_ipd;
      RDAD2_previous := RDAD2_ipd;
      RDAD1_previous := RDAD1_ipd;
      RDAD0_previous := RDAD0_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD7,
	GlitchData => RD7_GlitchData,
	OutSignalName => "RD7",
	OutTemp => RD7_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD7), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD7), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD7), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD7), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD7), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD7), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD7), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD7), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD7), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD7), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD7), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD7), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD7), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD7), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD7), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD7), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD7), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD7), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD7), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD7), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD7), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD7), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD7), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD7), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD7), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD6,
	GlitchData => RD6_GlitchData,
	OutSignalName => "RD6",
	OutTemp => RD6_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD6), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD6), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD6), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD6), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD6), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD6), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD6), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD6), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD6), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD6), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD6), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD6), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD6), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD6), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD6), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD6), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD6), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD6), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD6), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD6), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD6), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD6), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD6), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD6), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD6), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD5,
	GlitchData => RD5_GlitchData,
	OutSignalName => "RD5",
	OutTemp => RD5_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD5), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD5), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD5), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD5), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD5), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD5), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD5), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD5), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD5), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD5), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD5), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD5), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD5), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD5), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD5), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD5), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD5), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD5), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD5), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD5), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD5), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD5), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD5), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD5), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD5), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD4,
	GlitchData => RD4_GlitchData,
	OutSignalName => "RD4",
	OutTemp => RD4_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD4), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD4), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD4), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD4), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD4), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD4), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD4), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD4), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD4), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD4), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD4), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD4), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD4), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD4), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD4), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD4), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD4), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD4), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD4), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD4), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD4), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD4), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD4), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD4), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD4), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD3,
	GlitchData => RD3_GlitchData,
	OutSignalName => "RD3",
	OutTemp => RD3_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD2,
	GlitchData => RD2_GlitchData,
	OutSignalName => "RD2",
	OutTemp => RD2_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD1,
	GlitchData => RD1_GlitchData,
	OutSignalName => "RD1",
	OutTemp => RD1_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD0,
	GlitchData => RD0_GlitchData,
	OutSignalName => "RD0",
	OutTemp => RD0_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

  end process VITALBehavior;

end VITAL_ACT;
-----------------------------------------------------------------
--  Proxy Modeling, Inc. 
--
--  Actel RAM8FF VHDL behavioral model
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - Jan/22/96 - Initial Delivery
-- 1.1 - 12/6/96 by DNW - Modified SL_TO_INT.
-- 1.2 - 3/3/97 by DNW - WDx_delayed variables added.
-- 1.3 - 3/6/98 by DNW - Issue "unknown" msg. only if 0/1->X Xtion.
-- 1.4 - 5/27/98 by DNW - Initaialize _ipd signals to X instead of 0.
-- 
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity RAM8FF is
  GENERIC (
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD7      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD6      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD5      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD4      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD4_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC;
        RD6    : OUT STD_ULOGIC;
        RD5    : OUT STD_ULOGIC;
        RD4    : OUT STD_ULOGIC;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of RAM8FF : entity is TRUE;
  
end RAM8FF;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM8FF is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal WRAD4_ipd : std_ulogic := 'X';
  signal WRAD3_ipd : std_ulogic := 'X';
  signal WRAD2_ipd : std_ulogic := 'X';
  signal WRAD1_ipd : std_ulogic := 'X';
  signal WRAD0_ipd : std_ulogic := 'X';
  signal WD7_ipd : std_ulogic := 'X';
  signal WD6_ipd : std_ulogic := 'X';
  signal WD5_ipd : std_ulogic := 'X';
  signal WD4_ipd : std_ulogic := 'X';
  signal WD3_ipd : std_ulogic := 'X';
  signal WD2_ipd : std_ulogic := 'X';
  signal WD1_ipd : std_ulogic := 'X';
  signal WD0_ipd : std_ulogic := 'X';
  signal RDAD4_ipd : std_ulogic := 'X';
  signal RDAD3_ipd : std_ulogic := 'X';
  signal RDAD2_ipd : std_ulogic := 'X';
  signal RDAD1_ipd : std_ulogic := 'X';
  signal RDAD0_ipd : std_ulogic := 'X';
  signal BLKEN_ipd : std_ulogic := 'X';
  signal WEN_ipd : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal REN_ipd : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  type MEM is array(0 to 31) of std_ulogic_vector(7 downto 0);
   signal RAM_TMP : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (WRAD4_ipd, WRAD4, VitalExtendToFillDelay(tipd_WRAD4));
    VitalWireDelay (WRAD3_ipd, WRAD3, VitalExtendToFillDelay(tipd_WRAD3));
    VitalWireDelay (WRAD2_ipd, WRAD2, VitalExtendToFillDelay(tipd_WRAD2));
    VitalWireDelay (WRAD1_ipd, WRAD1, VitalExtendToFillDelay(tipd_WRAD1));
    VitalWireDelay (WRAD0_ipd, WRAD0, VitalExtendToFillDelay(tipd_WRAD0));
    VitalWireDelay (WD7_ipd, WD7, VitalExtendToFillDelay(tipd_WD7));
    VitalWireDelay (WD6_ipd, WD6, VitalExtendToFillDelay(tipd_WD6));
    VitalWireDelay (WD5_ipd, WD5, VitalExtendToFillDelay(tipd_WD5));
    VitalWireDelay (WD4_ipd, WD4, VitalExtendToFillDelay(tipd_WD4));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (RDAD4_ipd, RDAD4, VitalExtendToFillDelay(tipd_RDAD4));
    VitalWireDelay (RDAD3_ipd, RDAD3, VitalExtendToFillDelay(tipd_RDAD3));
    VitalWireDelay (RDAD2_ipd, RDAD2, VitalExtendToFillDelay(tipd_RDAD2));
    VitalWireDelay (RDAD1_ipd, RDAD1, VitalExtendToFillDelay(tipd_RDAD1));
    VitalWireDelay (RDAD0_ipd, RDAD0, VitalExtendToFillDelay(tipd_RDAD0));
    VitalWireDelay (BLKEN_ipd, BLKEN, VitalExtendToFillDelay(tipd_BLKEN));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (REN_ipd, REN, VitalExtendToFillDelay(tipd_REN));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (RDAD4_ipd, RDAD3_ipd, RDAD2_ipd, RDAD1_ipd, 
		RDAD0_ipd, REN_ipd, RCLK_ipd, WD7_ipd, WD6_ipd, WD5_ipd, 
		WD4_ipd, WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd, WRAD4_ipd, 
		WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, WEN_ipd, 
		BLKEN_ipd, BLKENS, WCLK_ipd)

     --  Read Timing Check Results
     variable Tviol_RDAD4_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD4_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD3_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD3_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD2_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD2_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD1_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD1_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD0_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD0_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_REN_RCLK_negedge : X01 := '0';
     variable TmDt_REN_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_WD7_WCLK_negedge : X01 := '0';
     variable TmDt_WD7_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD6_WCLK_negedge : X01 := '0';
     variable TmDt_WD6_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD5_WCLK_negedge : X01 := '0';
     variable TmDt_WD5_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD4_WCLK_negedge : X01 := '0';
     variable TmDt_WD4_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD3_WCLK_negedge : X01 := '0';
     variable TmDt_WD3_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_negedge : X01 := '0';
     variable TmDt_WD2_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_negedge : X01 := '0';
     variable TmDt_WD1_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_negedge : X01 := '0';
     variable TmDt_WD0_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD4_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD4_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD3_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD3_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD2_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD2_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD1_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD1_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD0_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD0_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_negedge : X01 := '0';
     variable TmDt_WEN_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_BLKEN_WCLK_negedge : X01 := '0';
     variable TmDt_BLKEN_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     --type SL_TO_INT is array(std_ulogic range <>) of integer;
     --constant INT :SL_TO_INT('U' to '-') := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     variable RD7_zd : std_ulogic;
     variable RD6_zd : std_ulogic;
     variable RD5_zd : std_ulogic;
     variable RD4_zd : std_ulogic;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD7_GlitchData : VitalGlitchDataType;
     variable RD6_GlitchData : VitalGlitchDataType;
     variable RD5_GlitchData : VitalGlitchDataType;
     variable RD4_GlitchData : VitalGlitchDataType;
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;
  
     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable WEN_delayed : std_ulogic := 'X';
     variable REN_delayed : std_ulogic := 'X';
     variable WEN_previous : std_ulogic := 'X';
     variable REN_previous : std_ulogic := 'X';
     variable BLKEN_delayed : std_ulogic := 'X';
     variable BLKEN_previous : std_ulogic := 'X';
     variable WD7_delayed : std_ulogic := 'X';
     variable WD6_delayed : std_ulogic := 'X';
     variable WD5_delayed : std_ulogic := 'X';
     variable WD4_delayed : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WRAD4_delayed : std_ulogic := 'X';
     variable WRAD3_delayed : std_ulogic := 'X';
     variable WRAD2_delayed : std_ulogic := 'X';
     variable WRAD1_delayed : std_ulogic := 'X';
     variable WRAD0_delayed : std_ulogic := 'X';
     variable WRAD4_previous : std_ulogic := 'X';
     variable WRAD3_previous : std_ulogic := 'X';
     variable WRAD2_previous : std_ulogic := 'X';
     variable WRAD1_previous : std_ulogic := 'X';
     variable WRAD0_previous : std_ulogic := 'X';
     variable RDAD4_delayed : std_ulogic := 'X';
     variable RDAD3_delayed : std_ulogic := 'X';
     variable RDAD2_delayed : std_ulogic := 'X';
     variable RDAD1_delayed : std_ulogic := 'X';
     variable RDAD0_delayed : std_ulogic := 'X';
     variable RDAD4_previous : std_ulogic := 'X';
     variable RDAD3_previous : std_ulogic := 'X';
     variable RDAD2_previous : std_ulogic := 'X';
     variable RDAD1_previous : std_ulogic := 'X';
     variable RDAD0_previous : std_ulogic := 'X';
  
  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RDAD high or low before RCLK falling
      --   Hold  RDAD high or low after RCLK falling

      VitalSetupHoldCheck ( Tviol_RDAD4_RCLK_negedge,
                            TmDt_RDAD4_RCLK_negedge,
                            RDAD4_ipd, "RDAD4",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD4_RCLK_noedge_negedge,
                            tsetup_RDAD4_RCLK_noedge_negedge,
                            thold_RDAD4_RCLK_noedge_negedge,
                            thold_RDAD4_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD3_RCLK_negedge,
                            TmDt_RDAD3_RCLK_negedge,
                            RDAD3_ipd, "RDAD3",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD3_RCLK_noedge_negedge,
                            tsetup_RDAD3_RCLK_noedge_negedge,
                            thold_RDAD3_RCLK_noedge_negedge,
                            thold_RDAD3_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD2_RCLK_negedge,
                            TmDt_RDAD2_RCLK_negedge,
                            RDAD2_ipd, "RDAD2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD2_RCLK_noedge_negedge,
                            tsetup_RDAD2_RCLK_noedge_negedge,
                            thold_RDAD2_RCLK_noedge_negedge,
                            thold_RDAD2_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD1_RCLK_negedge,
                            TmDt_RDAD1_RCLK_negedge,
                            RDAD1_ipd, "RDAD1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD1_RCLK_noedge_negedge,
                            tsetup_RDAD1_RCLK_noedge_negedge,
                            thold_RDAD1_RCLK_noedge_negedge,
                            thold_RDAD1_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD0_RCLK_negedge,
                            TmDt_RDAD0_RCLK_negedge,
                            RDAD0_ipd, "RDAD0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD0_RCLK_noedge_negedge,
                            tsetup_RDAD0_RCLK_noedge_negedge,
                            thold_RDAD0_RCLK_noedge_negedge,
                            thold_RDAD0_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup REN high before RCLK falling
      --   Hold  REN high after RCLK falling

      VitalSetupHoldCheck ( Tviol_REN_RCLK_negedge,
                            TmDt_REN_RCLK_negedge,
                            REN_ipd, "REN",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_REN_RCLK_noedge_negedge,
                            tsetup_REN_RCLK_noedge_negedge,
                            thold_REN_RCLK_noedge_negedge,
                            thold_REN_RCLK_noedge_negedge,
                            TimingCheckOn,
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup BLKEN high or low before WCLK falling
      --   Hold  BLKEN high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_BLKEN_WCLK_negedge,
                            TmDt_BLKEN_WCLK_negedge,
                            BLKEN_ipd, "BLKEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_BLKEN_WCLK_noedge_negedge,
                            tsetup_BLKEN_WCLK_noedge_negedge,
                            thold_BLKEN_WCLK_noedge_negedge,
                            thold_BLKEN_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WRAD high or low before WCLK falling
      --   Hold  WRAD high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_WRAD4_WCLK_negedge,
                            TmDt_WRAD4_WCLK_negedge,
                            WRAD4_ipd, "WRAD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD4_WCLK_noedge_negedge,
                            tsetup_WRAD4_WCLK_noedge_negedge,
                            thold_WRAD4_WCLK_noedge_negedge,
                            thold_WRAD4_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD3_WCLK_negedge,
                            TmDt_WRAD3_WCLK_negedge,
                            WRAD3_ipd, "WRAD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD3_WCLK_noedge_negedge,
                            tsetup_WRAD3_WCLK_noedge_negedge,
                            thold_WRAD3_WCLK_noedge_negedge,
                            thold_WRAD3_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD2_WCLK_negedge,
                            TmDt_WRAD2_WCLK_negedge,
                            WRAD2_ipd, "WRAD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD2_WCLK_noedge_negedge,
                            tsetup_WRAD2_WCLK_noedge_negedge,
                            thold_WRAD2_WCLK_noedge_negedge,
                            thold_WRAD2_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD1_WCLK_negedge,
                            TmDt_WRAD1_WCLK_negedge,
                            WRAD1_ipd, "WRAD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD1_WCLK_noedge_negedge,
                            tsetup_WRAD1_WCLK_noedge_negedge,
                            thold_WRAD1_WCLK_noedge_negedge,
                            thold_WRAD1_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD0_WCLK_negedge,
                            TmDt_WRAD0_WCLK_negedge,
                            WRAD0_ipd, "WRAD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD0_WCLK_noedge_negedge,
                            tsetup_WRAD0_WCLK_noedge_negedge,
                            thold_WRAD0_WCLK_noedge_negedge,
                            thold_WRAD0_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WD high or low before WCLK falling
      --   Hold  WD high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_WD7_WCLK_negedge,
                            TmDt_WD7_WCLK_negedge,
                            WD7_ipd, "WD7",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD7_WCLK_noedge_negedge,
                            tsetup_WD7_WCLK_noedge_negedge,
                            thold_WD7_WCLK_noedge_negedge,
                            thold_WD7_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD6_WCLK_negedge,
                            TmDt_WD6_WCLK_negedge,
                            WD6_ipd, "WD6",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD6_WCLK_noedge_negedge,
                            tsetup_WD6_WCLK_noedge_negedge,
                            thold_WD6_WCLK_noedge_negedge,
                            thold_WD6_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD5_WCLK_negedge,
                            TmDt_WD5_WCLK_negedge,
                            WD5_ipd, "WD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD5_WCLK_noedge_negedge,
                            tsetup_WD5_WCLK_noedge_negedge,
                            thold_WD5_WCLK_noedge_negedge,
                            thold_WD5_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD4_WCLK_negedge,
                            TmDt_WD4_WCLK_negedge,
                            WD4_ipd, "WD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD4_WCLK_noedge_negedge,
                            tsetup_WD4_WCLK_noedge_negedge,
                            thold_WD4_WCLK_noedge_negedge,
                            thold_WD4_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_negedge,
                            TmDt_WD3_WCLK_negedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_noedge_negedge,
                            tsetup_WD3_WCLK_noedge_negedge,
                            thold_WD3_WCLK_noedge_negedge,
                            thold_WD3_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_negedge,
                            TmDt_WD2_WCLK_negedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_noedge_negedge,
                            tsetup_WD2_WCLK_noedge_negedge,
                            thold_WD2_WCLK_noedge_negedge,
                            thold_WD2_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_negedge,
                            TmDt_WD1_WCLK_negedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_noedge_negedge,
                            tsetup_WD1_WCLK_noedge_negedge,
                            thold_WD1_WCLK_noedge_negedge,
                            thold_WD1_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_negedge,
                            TmDt_WD0_WCLK_negedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_noedge_negedge,
                            tsetup_WD0_WCLK_noedge_negedge,
                            thold_WD0_WCLK_noedge_negedge,
                            thold_WD0_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup WEN high before WCLK falling
      --   Hold  WEN high after WCLK falling

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_negedge,
                            TmDt_WEN_WCLK_negedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_noedge_negedge,
                            tsetup_WEN_WCLK_noedge_negedge,
                            thold_WEN_WCLK_noedge_negedge,
                            thold_WEN_WCLK_noedge_negedge,
                            (To_X01(BLKEN_ipd)=BLKENS),
                            '\',
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM8FF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
    
    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      -- Convert Write Address Signal to Integer
      WADDR := ((INT(WRAD4_delayed)*16)+(INT(WRAD3_delayed)*8)+(INT(WRAD2_delayed)*4)
		+(INT(WRAD1_delayed)*2)+(INT(WRAD0_delayed)));

      if (TO_X01(WCLK_ipd)='X') then
        if (TO_X01(WCLK_previous) /= 'X') then
	  assert false
	  report ": WCLK unknown"
	  severity Warning;
	end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='0')) then
	case TO_X01(WEN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (TO_X01(BLKEN_delayed) = 'X') then
              if (TO_X01(BLKEN_previous) /= 'X') then
	        assert false
	        report ": BLKEN unknown"
	        severity Warning;
	      end if;
	    elsif (TO_X01(BLKEN_delayed) = BLKENS) then
	      if (WADDR < 0) then
		if (TO_X01(WRAD4_delayed) = 'X') and (TO_X01(WRAD4_previous) /= 'X') then
		  assert false
		  report ": WRAD4 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD3_delayed) = 'X') and (TO_X01(WRAD3_previous) /= 'X') then
		  assert false
		  report ": WRAD3 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD2_delayed) = 'X') and (TO_X01(WRAD2_previous) /= 'X') then
		  assert false
		  report ": WRAD2 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD1_delayed) = 'X') and (TO_X01(WRAD1_previous) /= 'X') then
		  assert false
		  report ": WRAD1 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD0_delayed) = 'X') and (TO_X01(WRAD0_previous) /= 'X') then
		  assert false
		  report ": WRAD0 unknown"
		  severity Warning;
		end if;
	      else 
		RAM_TMP(WADDR) <= WD7_delayed & WD6_delayed & WD5_delayed & 
                                  WD4_delayed & WD3_delayed & WD2_delayed &
                                  WD1_delayed & WD0_delayed ; 
	      end if;
	    else
	      null;
	    end if;
	  when others =>
            if (TO_X01(WEN_previous) /= 'X') then
	      assert false
	      report ": WEN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      -- Convert Read Address Signal to Integer
      RADDR := ((INT(RDAD4_delayed)*16)+(INT(RDAD3_delayed)*8)+(INT(RDAD2_delayed)*4)
		+(INT(RDAD1_delayed)*2)+(INT(RDAD0_delayed)));

      if (TO_X01(RCLK_ipd) = 'X') then
	RD7_zd := 'X';
	RD6_zd := 'X';
	RD5_zd := 'X';
	RD4_zd := 'X';
	RD3_zd := 'X';
	RD2_zd := 'X';
	RD1_zd := 'X';
	RD0_zd := 'X';
	if (TO_X01(RCLK_previous) /= 'X') then
	  assert false
	  report ": RCLK unknown"
	  severity Warning;
	end if;
      elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '0')) then
	case TO_X01(REN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (RADDR < 0) then
	      RD7_zd := 'X';
	      RD6_zd := 'X';
	      RD5_zd := 'X';
	      RD4_zd := 'X';
	      RD3_zd := 'X';
	      RD2_zd := 'X';
	      RD1_zd := 'X';
	      RD0_zd := 'X';
	      if (TO_X01(RDAD4_delayed) = 'X') and (TO_X01(RDAD4_previous) /= 'X') then
		assert false
		report ": RDAD4 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD3_delayed) = 'X') and (TO_X01(RDAD3_previous) /= 'X') then
		assert false
		report ": RDAD3 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD2_delayed) = 'X') and (TO_X01(RDAD2_previous) /= 'X') then
		assert false
		report ": RDAD2 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD1_delayed) = 'X') and (TO_X01(RDAD1_previous) /= 'X') then
		assert false
		report ": RDAD1 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD0_delayed) = 'X') and (TO_X01(RDAD0_previous) /= 'X') then
		assert false
		report ": RDAD0 unknown"
		severity Warning;
	      end if;
	    else
	      RD7_zd := RAM_TMP(RADDR)(7);
	      RD6_zd := RAM_TMP(RADDR)(6);
	      RD5_zd := RAM_TMP(RADDR)(5);
	      RD4_zd := RAM_TMP(RADDR)(4);
	      RD3_zd := RAM_TMP(RADDR)(3);
	      RD2_zd := RAM_TMP(RADDR)(2);
	      RD1_zd := RAM_TMP(RADDR)(1);
	      RD0_zd := RAM_TMP(RADDR)(0);
	    end if;
	  when others =>
	    RD7_zd := 'X';
	    RD6_zd := 'X';
	    RD5_zd := 'X';
	    RD4_zd := 'X';
	    RD3_zd := 'X';
	    RD2_zd := 'X';
	    RD1_zd := 'X';
	    RD0_zd := 'X';
            if (TO_X01(REN_previous) /= 'X') then
	      assert false
	      report ": REN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;
      
      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      WEN_previous := WEN_delayed;
      REN_previous := REN_delayed;
      WEN_delayed := WEN_ipd;
      REN_delayed := REN_ipd;
      BLKEN_previous := BLKEN_delayed;
      BLKEN_delayed := BLKEN_ipd;
      WD7_delayed := WD7_ipd;
      WD6_delayed := WD6_ipd;
      WD5_delayed := WD5_ipd;
      WD4_delayed := WD4_ipd;
      WD3_delayed := WD3_ipd;
      WD2_delayed := WD2_ipd;
      WD1_delayed := WD1_ipd;
      WD0_delayed := WD0_ipd;
      WRAD4_previous := WRAD4_delayed;
      WRAD3_previous := WRAD3_delayed;
      WRAD2_previous := WRAD2_delayed;
      WRAD1_previous := WRAD1_delayed;
      WRAD0_previous := WRAD0_delayed;
      WRAD4_delayed := WRAD4_ipd;
      WRAD3_delayed := WRAD3_ipd;
      WRAD2_delayed := WRAD2_ipd;
      WRAD1_delayed := WRAD1_ipd;
      WRAD0_delayed := WRAD0_ipd;
      RDAD4_previous := RDAD4_delayed;
      RDAD3_previous := RDAD3_delayed;
      RDAD2_previous := RDAD2_delayed;
      RDAD1_previous := RDAD1_delayed;
      RDAD0_previous := RDAD0_delayed;
      RDAD4_delayed := RDAD4_ipd;
      RDAD3_delayed := RDAD3_ipd;
      RDAD2_delayed := RDAD2_ipd;
      RDAD1_delayed := RDAD1_ipd;
      RDAD0_delayed := RDAD0_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD7,
	GlitchData => RD7_GlitchData,
	OutSignalName => "RD7",
	OutTemp => RD7_zd,
	Paths => (0 => (RCLK_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RCLK_RD7), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD6,
	GlitchData => RD6_GlitchData,
	OutSignalName => "RD6",
	OutTemp => RD6_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD6), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD5,
	GlitchData => RD5_GlitchData,
	OutSignalName => "RD5",
	OutTemp => RD5_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD5), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD4,
	GlitchData => RD4_GlitchData,
	OutSignalName => "RD4",
	OutTemp => RD4_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD4), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD3,
	GlitchData => RD3_GlitchData,
	OutSignalName => "RD3",
	OutTemp => RD3_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD3), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD2,
	GlitchData => RD2_GlitchData,
	OutSignalName => "RD2",
	OutTemp => RD2_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD2), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD1,
	GlitchData => RD1_GlitchData,
	OutSignalName => "RD1",
	OutTemp => RD1_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD1), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD0,
	GlitchData => RD0_GlitchData,
	OutSignalName => "RD0",
	OutTemp => RD0_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD0), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

  end process VITALBehavior;

end VITAL_ACT;
-----------------------------------------------------------------
--  Proxy Modeling, Inc. 
--
--  Actel RAM8FR VHDL behavioral model
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - Jan/22/96 - Initial Delivery
-- 1.1 - 12/6/96 by DNW - Modified SL_TO_INT.
-- 1.2 - 3/3/97 by DNW - WDx_delayed variables added.
-- 1.3 - 3/6/98 by DNW - Issue "unknown" msg. only if 0/1->X Xtion.
-- 1.4 - 5/27/98 by DNW - Initaialize _ipd signals to X instead of 0.
-- 
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity RAM8FR is
  GENERIC (
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD7      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD6      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD5      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD4      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD4_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC;
        RD6    : OUT STD_ULOGIC;
        RD5    : OUT STD_ULOGIC;
        RD4    : OUT STD_ULOGIC;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of RAM8FR : entity is TRUE;
  
end RAM8FR;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM8FR is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal WRAD4_ipd : std_ulogic := 'X';
  signal WRAD3_ipd : std_ulogic := 'X';
  signal WRAD2_ipd : std_ulogic := 'X';
  signal WRAD1_ipd : std_ulogic := 'X';
  signal WRAD0_ipd : std_ulogic := 'X';
  signal WD7_ipd : std_ulogic := 'X';
  signal WD6_ipd : std_ulogic := 'X';
  signal WD5_ipd : std_ulogic := 'X';
  signal WD4_ipd : std_ulogic := 'X';
  signal WD3_ipd : std_ulogic := 'X';
  signal WD2_ipd : std_ulogic := 'X';
  signal WD1_ipd : std_ulogic := 'X';
  signal WD0_ipd : std_ulogic := 'X';
  signal RDAD4_ipd : std_ulogic := 'X';
  signal RDAD3_ipd : std_ulogic := 'X';
  signal RDAD2_ipd : std_ulogic := 'X';
  signal RDAD1_ipd : std_ulogic := 'X';
  signal RDAD0_ipd : std_ulogic := 'X';
  signal BLKEN_ipd : std_ulogic := 'X';
  signal WEN_ipd : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal REN_ipd : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  type MEM is array(0 to 31) of std_ulogic_vector(7 downto 0);
   signal RAM_TMP : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (WRAD4_ipd, WRAD4, VitalExtendToFillDelay(tipd_WRAD4));
    VitalWireDelay (WRAD3_ipd, WRAD3, VitalExtendToFillDelay(tipd_WRAD3));
    VitalWireDelay (WRAD2_ipd, WRAD2, VitalExtendToFillDelay(tipd_WRAD2));
    VitalWireDelay (WRAD1_ipd, WRAD1, VitalExtendToFillDelay(tipd_WRAD1));
    VitalWireDelay (WRAD0_ipd, WRAD0, VitalExtendToFillDelay(tipd_WRAD0));
    VitalWireDelay (WD7_ipd, WD7, VitalExtendToFillDelay(tipd_WD7));
    VitalWireDelay (WD6_ipd, WD6, VitalExtendToFillDelay(tipd_WD6));
    VitalWireDelay (WD5_ipd, WD5, VitalExtendToFillDelay(tipd_WD5));
    VitalWireDelay (WD4_ipd, WD4, VitalExtendToFillDelay(tipd_WD4));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (RDAD4_ipd, RDAD4, VitalExtendToFillDelay(tipd_RDAD4));
    VitalWireDelay (RDAD3_ipd, RDAD3, VitalExtendToFillDelay(tipd_RDAD3));
    VitalWireDelay (RDAD2_ipd, RDAD2, VitalExtendToFillDelay(tipd_RDAD2));
    VitalWireDelay (RDAD1_ipd, RDAD1, VitalExtendToFillDelay(tipd_RDAD1));
    VitalWireDelay (RDAD0_ipd, RDAD0, VitalExtendToFillDelay(tipd_RDAD0));
    VitalWireDelay (BLKEN_ipd, BLKEN, VitalExtendToFillDelay(tipd_BLKEN));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (REN_ipd, REN, VitalExtendToFillDelay(tipd_REN));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (RDAD4_ipd, RDAD3_ipd, RDAD2_ipd, RDAD1_ipd, 
		RDAD0_ipd, REN_ipd, RCLK_ipd, WD7_ipd, WD6_ipd, WD5_ipd, 
		WD4_ipd, WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd, WRAD4_ipd, 
		WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, WEN_ipd, 
		BLKEN_ipd, BLKENS, WCLK_ipd)

     --  Read Timing Check Results
     variable Tviol_RDAD4_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD4_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD3_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD2_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD1_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD0_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_REN_RCLK_posedge : X01 := '0';
     variable TmDt_REN_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_WD7_WCLK_negedge : X01 := '0';
     variable TmDt_WD7_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD6_WCLK_negedge : X01 := '0';
     variable TmDt_WD6_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD5_WCLK_negedge : X01 := '0';
     variable TmDt_WD5_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD4_WCLK_negedge : X01 := '0';
     variable TmDt_WD4_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD3_WCLK_negedge : X01 := '0';
     variable TmDt_WD3_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_negedge : X01 := '0';
     variable TmDt_WD2_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_negedge : X01 := '0';
     variable TmDt_WD1_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_negedge : X01 := '0';
     variable TmDt_WD0_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD4_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD4_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD3_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD3_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD2_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD2_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD1_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD1_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD0_WCLK_negedge : X01 := '0';
     variable TmDt_WRAD0_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_negedge : X01 := '0';
     variable TmDt_WEN_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_BLKEN_WCLK_negedge : X01 := '0';
     variable TmDt_BLKEN_WCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     --type SL_TO_INT is array(std_ulogic range <>) of integer;
     --constant INT :SL_TO_INT('U' to '-') := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     variable RD7_zd : std_ulogic;
     variable RD6_zd : std_ulogic;
     variable RD5_zd : std_ulogic;
     variable RD4_zd : std_ulogic;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD7_GlitchData : VitalGlitchDataType;
     variable RD6_GlitchData : VitalGlitchDataType;
     variable RD5_GlitchData : VitalGlitchDataType;
     variable RD4_GlitchData : VitalGlitchDataType;
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;
  
     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable WEN_delayed : std_ulogic := 'X';
     variable REN_delayed : std_ulogic := 'X';
     variable WEN_previous : std_ulogic := 'X';
     variable REN_previous : std_ulogic := 'X';
     variable BLKEN_delayed : std_ulogic := 'X';
     variable BLKEN_previous : std_ulogic := 'X';
     variable WD7_delayed : std_ulogic := 'X';
     variable WD6_delayed : std_ulogic := 'X';
     variable WD5_delayed : std_ulogic := 'X';
     variable WD4_delayed : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WRAD4_delayed : std_ulogic := 'X';
     variable WRAD3_delayed : std_ulogic := 'X';
     variable WRAD2_delayed : std_ulogic := 'X';
     variable WRAD1_delayed : std_ulogic := 'X';
     variable WRAD0_delayed : std_ulogic := 'X';
     variable WRAD4_previous : std_ulogic := 'X';
     variable WRAD3_previous : std_ulogic := 'X';
     variable WRAD2_previous : std_ulogic := 'X';
     variable WRAD1_previous : std_ulogic := 'X';
     variable WRAD0_previous : std_ulogic := 'X';
     variable RDAD4_delayed : std_ulogic := 'X';
     variable RDAD3_delayed : std_ulogic := 'X';
     variable RDAD2_delayed : std_ulogic := 'X';
     variable RDAD1_delayed : std_ulogic := 'X';
     variable RDAD0_delayed : std_ulogic := 'X';
     variable RDAD4_previous : std_ulogic := 'X';
     variable RDAD3_previous : std_ulogic := 'X';
     variable RDAD2_previous : std_ulogic := 'X';
     variable RDAD1_previous : std_ulogic := 'X';
     variable RDAD0_previous : std_ulogic := 'X';
  
  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RDAD high or low before RCLK rising
      --   Hold  RDAD high or low after RCLK rising

      VitalSetupHoldCheck ( Tviol_RDAD4_RCLK_posedge,
                            TmDt_RDAD4_RCLK_posedge,
                            RDAD4_ipd, "RDAD4",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD4_RCLK_noedge_posedge,
                            tsetup_RDAD4_RCLK_noedge_posedge,
                            thold_RDAD4_RCLK_noedge_posedge,
                            thold_RDAD4_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD3_RCLK_posedge,
                            TmDt_RDAD3_RCLK_posedge,
                            RDAD3_ipd, "RDAD3",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD3_RCLK_noedge_posedge,
                            tsetup_RDAD3_RCLK_noedge_posedge,
                            thold_RDAD3_RCLK_noedge_posedge,
                            thold_RDAD3_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD2_RCLK_posedge,
                            TmDt_RDAD2_RCLK_posedge,
                            RDAD2_ipd, "RDAD2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD2_RCLK_noedge_posedge,
                            tsetup_RDAD2_RCLK_noedge_posedge,
                            thold_RDAD2_RCLK_noedge_posedge,
                            thold_RDAD2_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD1_RCLK_posedge,
                            TmDt_RDAD1_RCLK_posedge,
                            RDAD1_ipd, "RDAD1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD1_RCLK_noedge_posedge,
                            tsetup_RDAD1_RCLK_noedge_posedge,
                            thold_RDAD1_RCLK_noedge_posedge,
                            thold_RDAD1_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD0_RCLK_posedge,
                            TmDt_RDAD0_RCLK_posedge,
                            RDAD0_ipd, "RDAD0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD0_RCLK_noedge_posedge,
                            tsetup_RDAD0_RCLK_noedge_posedge,
                            thold_RDAD0_RCLK_noedge_posedge,
                            thold_RDAD0_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup REN high before RCLK rising
      --   Hold  REN high after RCLK rising

      VitalSetupHoldCheck ( Tviol_REN_RCLK_posedge,
                            TmDt_REN_RCLK_posedge,
                            REN_ipd, "REN",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_REN_RCLK_noedge_posedge,
                            tsetup_REN_RCLK_noedge_posedge,
                            thold_REN_RCLK_noedge_posedge,
                            thold_REN_RCLK_noedge_posedge,
                            TimingCheckOn,
                            '/',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup BLKEN high or low before WCLK falling
      --   Hold  BLKEN high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_BLKEN_WCLK_negedge,
                            TmDt_BLKEN_WCLK_negedge,
                            BLKEN_ipd, "BLKEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_BLKEN_WCLK_noedge_negedge,
                            tsetup_BLKEN_WCLK_noedge_negedge,
                            thold_BLKEN_WCLK_noedge_negedge,
                            thold_BLKEN_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WRAD high or low before WCLK falling
      --   Hold  WRAD high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_WRAD4_WCLK_negedge,
                            TmDt_WRAD4_WCLK_negedge,
                            WRAD4_ipd, "WRAD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD4_WCLK_noedge_negedge,
                            tsetup_WRAD4_WCLK_noedge_negedge,
                            thold_WRAD4_WCLK_noedge_negedge,
                            thold_WRAD4_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD3_WCLK_negedge,
                            TmDt_WRAD3_WCLK_negedge,
                            WRAD3_ipd, "WRAD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD3_WCLK_noedge_negedge,
                            tsetup_WRAD3_WCLK_noedge_negedge,
                            thold_WRAD3_WCLK_noedge_negedge,
                            thold_WRAD3_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD2_WCLK_negedge,
                            TmDt_WRAD2_WCLK_negedge,
                            WRAD2_ipd, "WRAD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD2_WCLK_noedge_negedge,
                            tsetup_WRAD2_WCLK_noedge_negedge,
                            thold_WRAD2_WCLK_noedge_negedge,
                            thold_WRAD2_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD1_WCLK_negedge,
                            TmDt_WRAD1_WCLK_negedge,
                            WRAD1_ipd, "WRAD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD1_WCLK_noedge_negedge,
                            tsetup_WRAD1_WCLK_noedge_negedge,
                            thold_WRAD1_WCLK_noedge_negedge,
                            thold_WRAD1_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD0_WCLK_negedge,
                            TmDt_WRAD0_WCLK_negedge,
                            WRAD0_ipd, "WRAD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD0_WCLK_noedge_negedge,
                            tsetup_WRAD0_WCLK_noedge_negedge,
                            thold_WRAD0_WCLK_noedge_negedge,
                            thold_WRAD0_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WD high or low before WCLK falling
      --   Hold  WD high or low before WCLK falling

      VitalSetupHoldCheck ( Tviol_WD7_WCLK_negedge,
                            TmDt_WD7_WCLK_negedge,
                            WD7_ipd, "WD7",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD7_WCLK_noedge_negedge,
                            tsetup_WD7_WCLK_noedge_negedge,
                            thold_WD7_WCLK_noedge_negedge,
                            thold_WD7_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD6_WCLK_negedge,
                            TmDt_WD6_WCLK_negedge,
                            WD6_ipd, "WD6",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD6_WCLK_noedge_negedge,
                            tsetup_WD6_WCLK_noedge_negedge,
                            thold_WD6_WCLK_noedge_negedge,
                            thold_WD6_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD5_WCLK_negedge,
                            TmDt_WD5_WCLK_negedge,
                            WD5_ipd, "WD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD5_WCLK_noedge_negedge,
                            tsetup_WD5_WCLK_noedge_negedge,
                            thold_WD5_WCLK_noedge_negedge,
                            thold_WD5_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD4_WCLK_negedge,
                            TmDt_WD4_WCLK_negedge,
                            WD4_ipd, "WD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD4_WCLK_noedge_negedge,
                            tsetup_WD4_WCLK_noedge_negedge,
                            thold_WD4_WCLK_noedge_negedge,
                            thold_WD4_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_negedge,
                            TmDt_WD3_WCLK_negedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_noedge_negedge,
                            tsetup_WD3_WCLK_noedge_negedge,
                            thold_WD3_WCLK_noedge_negedge,
                            thold_WD3_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_negedge,
                            TmDt_WD2_WCLK_negedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_noedge_negedge,
                            tsetup_WD2_WCLK_noedge_negedge,
                            thold_WD2_WCLK_noedge_negedge,
                            thold_WD2_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_negedge,
                            TmDt_WD1_WCLK_negedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_noedge_negedge,
                            tsetup_WD1_WCLK_noedge_negedge,
                            thold_WD1_WCLK_noedge_negedge,
                            thold_WD1_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_negedge,
                            TmDt_WD0_WCLK_negedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_noedge_negedge,
                            tsetup_WD0_WCLK_noedge_negedge,
                            thold_WD0_WCLK_noedge_negedge,
                            thold_WD0_WCLK_noedge_negedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup WEN high before WCLK falling
      --   Hold  WEN high after WCLK falling

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_negedge,
                            TmDt_WEN_WCLK_negedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_noedge_negedge,
                            tsetup_WEN_WCLK_noedge_negedge,
                            thold_WEN_WCLK_noedge_negedge,
                            thold_WEN_WCLK_noedge_negedge,
                            (To_X01(BLKEN_ipd)=BLKENS),
                            '\',
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM8FR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
    
    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      -- Convert Write Address Signal to Integer
      WADDR := ((INT(WRAD4_delayed)*16)+(INT(WRAD3_delayed)*8)+(INT(WRAD2_delayed)*4)
		+(INT(WRAD1_delayed)*2)+(INT(WRAD0_delayed)));

      if (TO_X01(WCLK_ipd)='X') then
        if (TO_X01(WCLK_previous) /= 'X') then
	  assert false
	  report ": WCLK unknown"
	  severity Warning;
	end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='0')) then
	case TO_X01(WEN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (TO_X01(BLKEN_delayed) = 'X') then
              if (TO_X01(BLKEN_previous) /= 'X') then
	        assert false
	        report ": BLKEN unknown"
	        severity Warning;
	      end if;
	    elsif (TO_X01(BLKEN_delayed) = BLKENS) then
	      if (WADDR < 0) then
		if (TO_X01(WRAD4_delayed) = 'X') and (TO_X01(WRAD4_previous) /= 'X') then
		  assert false
		  report ": WRAD4 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD3_delayed) = 'X') and (TO_X01(WRAD3_previous) /= 'X') then
		  assert false
		  report ": WRAD3 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD2_delayed) = 'X') and (TO_X01(WRAD2_previous) /= 'X') then
		  assert false
		  report ": WRAD2 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD1_delayed) = 'X') and (TO_X01(WRAD1_previous) /= 'X') then
		  assert false
		  report ": WRAD1 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD0_delayed) = 'X') and (TO_X01(WRAD0_previous) /= 'X') then
		  assert false
		  report ": WRAD0 unknown"
		  severity Warning;
		end if;
	      else 
		RAM_TMP(WADDR) <= WD7_delayed & WD6_delayed & WD5_delayed & 
                                  WD4_delayed & WD3_delayed & WD2_delayed &
                                  WD1_delayed & WD0_delayed ; 
	      end if;
	    else
	      null;
	    end if;
	  when others =>
            if (TO_X01(WEN_previous) /= 'X') then
	      assert false
	      report ": WEN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      -- Convert Read Address Signal to Integer
      RADDR := ((INT(RDAD4_delayed)*16)+(INT(RDAD3_delayed)*8)+(INT(RDAD2_delayed)*4)
		+(INT(RDAD1_delayed)*2)+(INT(RDAD0_delayed)));

      if (TO_X01(RCLK_ipd) = 'X') then
	RD7_zd := 'X';
	RD6_zd := 'X';
	RD5_zd := 'X';
	RD4_zd := 'X';
	RD3_zd := 'X';
	RD2_zd := 'X';
	RD1_zd := 'X';
	RD0_zd := 'X';
	if (TO_X01(RCLK_previous) /= 'X') then
	  assert false
	  report ": RCLK unknown"
	  severity Warning;
	end if;
      elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1')) then
	case TO_X01(REN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (RADDR < 0) then
	      RD7_zd := 'X';
	      RD6_zd := 'X';
	      RD5_zd := 'X';
	      RD4_zd := 'X';
	      RD3_zd := 'X';
	      RD2_zd := 'X';
	      RD1_zd := 'X';
	      RD0_zd := 'X';
	      if (TO_X01(RDAD4_delayed) = 'X') and (TO_X01(RDAD4_previous) /= 'X') then
		assert false
		report ": RDAD4 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD3_delayed) = 'X') and (TO_X01(RDAD3_previous) /= 'X') then
		assert false
		report ": RDAD3 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD2_delayed) = 'X') and (TO_X01(RDAD2_previous) /= 'X') then
		assert false
		report ": RDAD2 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD1_delayed) = 'X') and (TO_X01(RDAD1_previous) /= 'X') then
		assert false
		report ": RDAD1 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD0_delayed) = 'X') and (TO_X01(RDAD0_previous) /= 'X') then
		assert false
		report ": RDAD0 unknown"
		severity Warning;
	      end if;
	    else
	      RD7_zd := RAM_TMP(RADDR)(7);
	      RD6_zd := RAM_TMP(RADDR)(6);
	      RD5_zd := RAM_TMP(RADDR)(5);
	      RD4_zd := RAM_TMP(RADDR)(4);
	      RD3_zd := RAM_TMP(RADDR)(3);
	      RD2_zd := RAM_TMP(RADDR)(2);
	      RD1_zd := RAM_TMP(RADDR)(1);
	      RD0_zd := RAM_TMP(RADDR)(0);
	    end if;
	  when others =>
	    RD7_zd := 'X';
	    RD6_zd := 'X';
	    RD5_zd := 'X';
	    RD4_zd := 'X';
	    RD3_zd := 'X';
	    RD2_zd := 'X';
	    RD1_zd := 'X';
	    RD0_zd := 'X';
            if (TO_X01(REN_previous) /= 'X') then
	      assert false
	      report ": REN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;
      
      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      WEN_previous := WEN_delayed;
      REN_previous := REN_delayed;
      WEN_delayed := WEN_ipd;
      REN_delayed := REN_ipd;
      BLKEN_previous := BLKEN_delayed;
      BLKEN_delayed := BLKEN_ipd;
      WD7_delayed := WD7_ipd;
      WD6_delayed := WD6_ipd;
      WD5_delayed := WD5_ipd;
      WD4_delayed := WD4_ipd;
      WD3_delayed := WD3_ipd;
      WD2_delayed := WD2_ipd;
      WD1_delayed := WD1_ipd;
      WD0_delayed := WD0_ipd;
      WRAD4_previous := WRAD4_delayed;
      WRAD3_previous := WRAD3_delayed;
      WRAD2_previous := WRAD2_delayed;
      WRAD1_previous := WRAD1_delayed;
      WRAD0_previous := WRAD0_delayed;
      WRAD4_delayed := WRAD4_ipd;
      WRAD3_delayed := WRAD3_ipd;
      WRAD2_delayed := WRAD2_ipd;
      WRAD1_delayed := WRAD1_ipd;
      WRAD0_delayed := WRAD0_ipd;
      RDAD4_previous := RDAD4_delayed;
      RDAD3_previous := RDAD3_delayed;
      RDAD2_previous := RDAD2_delayed;
      RDAD1_previous := RDAD1_delayed;
      RDAD0_previous := RDAD0_delayed;
      RDAD4_delayed := RDAD4_ipd;
      RDAD3_delayed := RDAD3_ipd;
      RDAD2_delayed := RDAD2_ipd;
      RDAD1_delayed := RDAD1_ipd;
      RDAD0_delayed := RDAD0_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD7,
	GlitchData => RD7_GlitchData,
	OutSignalName => "RD7",
	OutTemp => RD7_zd,
	Paths => (0 => (RCLK_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RCLK_RD7), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD6,
	GlitchData => RD6_GlitchData,
	OutSignalName => "RD6",
	OutTemp => RD6_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD6), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD5,
	GlitchData => RD5_GlitchData,
	OutSignalName => "RD5",
	OutTemp => RD5_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD5), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD4,
	GlitchData => RD4_GlitchData,
	OutSignalName => "RD4",
	OutTemp => RD4_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD4), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD3,
	GlitchData => RD3_GlitchData,
	OutSignalName => "RD3",
	OutTemp => RD3_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD3), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD2,
	GlitchData => RD2_GlitchData,
	OutSignalName => "RD2",
	OutTemp => RD2_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD2), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD1,
	GlitchData => RD1_GlitchData,
	OutSignalName => "RD1",
	OutTemp => RD1_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD1), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD0,
	GlitchData => RD0_GlitchData,
	OutSignalName => "RD0",
	OutTemp => RD0_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD0), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

  end process VITALBehavior;

end VITAL_ACT;
-----------------------------------------------------------------
--  Proxy Modeling, Inc. 
--
--  Actel RAM8RA VHDL behavioral model
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - Jan/22/96 - Initial Delivery
-- 1.1 - 12/6/96 by DNW - Modified SL_TO_INT.
-- 1.2 - 3/3/97 by DNW - WDx_delayed variables added.
-- 1.3 - 3/6/98 by DNW - Issue "unknown" msg. only if 0/1->X Xtion.
-- 1.4 - 5/27/98 by DNW - Initaialize _ipd signals to X instead of 0.
-- 
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity RAM8RA is
  GENERIC (
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD7      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD6      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD5      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD4      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RDAD4_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD4_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD3_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD2_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD1_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RDAD0_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_WRAD4_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC;
        RD6    : OUT STD_ULOGIC;
        RD5    : OUT STD_ULOGIC;
        RD4    : OUT STD_ULOGIC;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of RAM8RA : entity is TRUE;
  
end RAM8RA;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM8RA is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal WRAD4_ipd : std_ulogic := 'X';
  signal WRAD3_ipd : std_ulogic := 'X';
  signal WRAD2_ipd : std_ulogic := 'X';
  signal WRAD1_ipd : std_ulogic := 'X';
  signal WRAD0_ipd : std_ulogic := 'X';
  signal WD7_ipd : std_ulogic := 'X';
  signal WD6_ipd : std_ulogic := 'X';
  signal WD5_ipd : std_ulogic := 'X';
  signal WD4_ipd : std_ulogic := 'X';
  signal WD3_ipd : std_ulogic := 'X';
  signal WD2_ipd : std_ulogic := 'X';
  signal WD1_ipd : std_ulogic := 'X';
  signal WD0_ipd : std_ulogic := 'X';
  signal RDAD4_ipd : std_ulogic := 'X';
  signal RDAD3_ipd : std_ulogic := 'X';
  signal RDAD2_ipd : std_ulogic := 'X';
  signal RDAD1_ipd : std_ulogic := 'X';
  signal RDAD0_ipd : std_ulogic := 'X';
  signal BLKEN_ipd : std_ulogic := 'X';
  signal WEN_ipd : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  type MEM is array(0 to 31) of std_ulogic_vector(7 downto 0);
   signal RAM_TMP : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (WRAD4_ipd, WRAD4, VitalExtendToFillDelay(tipd_WRAD4));
    VitalWireDelay (WRAD3_ipd, WRAD3, VitalExtendToFillDelay(tipd_WRAD3));
    VitalWireDelay (WRAD2_ipd, WRAD2, VitalExtendToFillDelay(tipd_WRAD2));
    VitalWireDelay (WRAD1_ipd, WRAD1, VitalExtendToFillDelay(tipd_WRAD1));
    VitalWireDelay (WRAD0_ipd, WRAD0, VitalExtendToFillDelay(tipd_WRAD0));
    VitalWireDelay (WD7_ipd, WD7, VitalExtendToFillDelay(tipd_WD7));
    VitalWireDelay (WD6_ipd, WD6, VitalExtendToFillDelay(tipd_WD6));
    VitalWireDelay (WD5_ipd, WD5, VitalExtendToFillDelay(tipd_WD5));
    VitalWireDelay (WD4_ipd, WD4, VitalExtendToFillDelay(tipd_WD4));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (RDAD4_ipd, RDAD4, VitalExtendToFillDelay(tipd_RDAD4));
    VitalWireDelay (RDAD3_ipd, RDAD3, VitalExtendToFillDelay(tipd_RDAD3));
    VitalWireDelay (RDAD2_ipd, RDAD2, VitalExtendToFillDelay(tipd_RDAD2));
    VitalWireDelay (RDAD1_ipd, RDAD1, VitalExtendToFillDelay(tipd_RDAD1));
    VitalWireDelay (RDAD0_ipd, RDAD0, VitalExtendToFillDelay(tipd_RDAD0));
    VitalWireDelay (BLKEN_ipd, BLKEN, VitalExtendToFillDelay(tipd_BLKEN));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (RDAD4_ipd, RDAD3_ipd, RDAD2_ipd, RDAD1_ipd, 
		RDAD0_ipd, WD7_ipd, WD6_ipd, WD5_ipd, 
		WD4_ipd, WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd, WRAD4_ipd, 
		WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, WEN_ipd, 
		BLKEN_ipd, BLKENS, WCLK_ipd, RAM_TMP)

     --  Write Timing Check Results
     variable Tviol_WD7_WCLK_posedge : X01 := '0';
     variable TmDt_WD7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD6_WCLK_posedge : X01 := '0';
     variable TmDt_WD6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD5_WCLK_posedge : X01 := '0';
     variable TmDt_WD5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD4_WCLK_posedge : X01 := '0';
     variable TmDt_WD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD3_WCLK_posedge : X01 := '0';
     variable TmDt_WD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_posedge : X01 := '0';
     variable TmDt_WD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_posedge : X01 := '0';
     variable TmDt_WD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_posedge : X01 := '0';
     variable TmDt_WD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD4_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD3_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD2_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD1_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD0_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_posedge : X01 := '0';
     variable TmDt_WEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_BLKEN_WCLK_posedge : X01 := '0';
     variable TmDt_BLKEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     --type SL_TO_INT is array(std_ulogic range <>) of integer;
     --constant INT :SL_TO_INT('U' to '-') := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     variable RD7_zd : std_ulogic;
     variable RD6_zd : std_ulogic;
     variable RD5_zd : std_ulogic;
     variable RD4_zd : std_ulogic;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD7_GlitchData : VitalGlitchDataType;
     variable RD6_GlitchData : VitalGlitchDataType;
     variable RD5_GlitchData : VitalGlitchDataType;
     variable RD4_GlitchData : VitalGlitchDataType;
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;
  
     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable WEN_delayed : std_ulogic := 'X';
     variable WEN_previous : std_ulogic := 'X';
     variable BLKEN_delayed : std_ulogic := 'X';
     variable BLKEN_previous : std_ulogic := 'X';
     variable WD7_delayed : std_ulogic := 'X';
     variable WD6_delayed : std_ulogic := 'X';
     variable WD5_delayed : std_ulogic := 'X';
     variable WD4_delayed : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WRAD4_delayed : std_ulogic := 'X';
     variable WRAD3_delayed : std_ulogic := 'X';
     variable WRAD2_delayed : std_ulogic := 'X';
     variable WRAD1_delayed : std_ulogic := 'X';
     variable WRAD0_delayed : std_ulogic := 'X';
     variable WRAD4_previous : std_ulogic := 'X';
     variable WRAD3_previous : std_ulogic := 'X';
     variable WRAD2_previous : std_ulogic := 'X';
     variable WRAD1_previous : std_ulogic := 'X';
     variable WRAD0_previous : std_ulogic := 'X';
     variable RDAD4_previous : std_ulogic := 'X';
     variable RDAD3_previous : std_ulogic := 'X';
     variable RDAD2_previous : std_ulogic := 'X';
     variable RDAD1_previous : std_ulogic := 'X';
     variable RDAD0_previous : std_ulogic := 'X';
  
  begin  --  process VITALBehavior 

    if (TimingCheckOn) then

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup BLKEN high or low before WCLK rising
      --   Hold  BLKEN high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_BLKEN_WCLK_posedge,
                            TmDt_BLKEN_WCLK_posedge,
                            BLKEN_ipd, "BLKEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_BLKEN_WCLK_noedge_posedge,
                            tsetup_BLKEN_WCLK_noedge_posedge,
                            thold_BLKEN_WCLK_noedge_posedge,
                            thold_BLKEN_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WRAD high or low before WCLK rising
      --   Hold  WRAD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WRAD4_WCLK_posedge,
                            TmDt_WRAD4_WCLK_posedge,
                            WRAD4_ipd, "WRAD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD4_WCLK_noedge_posedge,
                            tsetup_WRAD4_WCLK_noedge_posedge,
                            thold_WRAD4_WCLK_noedge_posedge,
                            thold_WRAD4_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD3_WCLK_posedge,
                            TmDt_WRAD3_WCLK_posedge,
                            WRAD3_ipd, "WRAD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD3_WCLK_noedge_posedge,
                            tsetup_WRAD3_WCLK_noedge_posedge,
                            thold_WRAD3_WCLK_noedge_posedge,
                            thold_WRAD3_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD2_WCLK_posedge,
                            TmDt_WRAD2_WCLK_posedge,
                            WRAD2_ipd, "WRAD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD2_WCLK_noedge_posedge,
                            tsetup_WRAD2_WCLK_noedge_posedge,
                            thold_WRAD2_WCLK_noedge_posedge,
                            thold_WRAD2_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD1_WCLK_posedge,
                            TmDt_WRAD1_WCLK_posedge,
                            WRAD1_ipd, "WRAD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD1_WCLK_noedge_posedge,
                            tsetup_WRAD1_WCLK_noedge_posedge,
                            thold_WRAD1_WCLK_noedge_posedge,
                            thold_WRAD1_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD0_WCLK_posedge,
                            TmDt_WRAD0_WCLK_posedge,
                            WRAD0_ipd, "WRAD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD0_WCLK_noedge_posedge,
                            tsetup_WRAD0_WCLK_noedge_posedge,
                            thold_WRAD0_WCLK_noedge_posedge,
                            thold_WRAD0_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WD high or low before WCLK rising
      --   Hold  WD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WD7_WCLK_posedge,
                            TmDt_WD7_WCLK_posedge,
                            WD7_ipd, "WD7",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD7_WCLK_noedge_posedge,
                            tsetup_WD7_WCLK_noedge_posedge,
                            thold_WD7_WCLK_noedge_posedge,
                            thold_WD7_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD6_WCLK_posedge,
                            TmDt_WD6_WCLK_posedge,
                            WD6_ipd, "WD6",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD6_WCLK_noedge_posedge,
                            tsetup_WD6_WCLK_noedge_posedge,
                            thold_WD6_WCLK_noedge_posedge,
                            thold_WD6_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD5_WCLK_posedge,
                            TmDt_WD5_WCLK_posedge,
                            WD5_ipd, "WD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD5_WCLK_noedge_posedge,
                            tsetup_WD5_WCLK_noedge_posedge,
                            thold_WD5_WCLK_noedge_posedge,
                            thold_WD5_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD4_WCLK_posedge,
                            TmDt_WD4_WCLK_posedge,
                            WD4_ipd, "WD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD4_WCLK_noedge_posedge,
                            tsetup_WD4_WCLK_noedge_posedge,
                            thold_WD4_WCLK_noedge_posedge,
                            thold_WD4_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_posedge,
                            TmDt_WD3_WCLK_posedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_noedge_posedge,
                            tsetup_WD3_WCLK_noedge_posedge,
                            thold_WD3_WCLK_noedge_posedge,
                            thold_WD3_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_posedge,
                            TmDt_WD2_WCLK_posedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_noedge_posedge,
                            tsetup_WD2_WCLK_noedge_posedge,
                            thold_WD2_WCLK_noedge_posedge,
                            thold_WD2_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_posedge,
                            TmDt_WD1_WCLK_posedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_noedge_posedge,
                            tsetup_WD1_WCLK_noedge_posedge,
                            thold_WD1_WCLK_noedge_posedge,
                            thold_WD1_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_posedge,
                            TmDt_WD0_WCLK_posedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_noedge_posedge,
                            tsetup_WD0_WCLK_noedge_posedge,
                            thold_WD0_WCLK_noedge_posedge,
                            thold_WD0_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup WEN high before WCLK rising
      --   Hold  WEN high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_posedge,
                            TmDt_WEN_WCLK_posedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_noedge_posedge,
                            tsetup_WEN_WCLK_noedge_posedge,
                            thold_WEN_WCLK_noedge_posedge,
                            thold_WEN_WCLK_noedge_posedge,
                            (To_X01(BLKEN_ipd)=BLKENS),
                            '/',
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM8RA",
                            TRUE,
                            TRUE,
                            ERROR
                            );
    
    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      -- Convert Write Address Signal to Integer
      WADDR := ((INT(WRAD4_delayed)*16)+(INT(WRAD3_delayed)*8)+(INT(WRAD2_delayed)*4)
		+(INT(WRAD1_delayed)*2)+(INT(WRAD0_delayed)));

      if (TO_X01(WCLK_ipd)='X') then
        if (TO_X01(WCLK_previous) /= 'X') then
	  assert false
	  report ": WCLK unknown"
	  severity Warning;
	end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	case TO_X01(WEN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (TO_X01(BLKEN_delayed) = 'X') then
              if (TO_X01(BLKEN_previous) /= 'X') then
	        assert false
	        report ": BLKEN unknown"
	        severity Warning;
	      end if;
	    elsif (TO_X01(BLKEN_delayed) = BLKENS) then
	      if (WADDR < 0) then
		if (TO_X01(WRAD4_delayed) = 'X') and (TO_X01(WRAD4_previous) /= 'X') then
		  assert false
		  report ": WRAD4 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD3_delayed) = 'X') and (TO_X01(WRAD3_previous) /= 'X') then
		  assert false
		  report ": WRAD3 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD2_delayed) = 'X') and (TO_X01(WRAD2_previous) /= 'X') then
		  assert false
		  report ": WRAD2 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD1_delayed) = 'X') and (TO_X01(WRAD1_previous) /= 'X') then
		  assert false
		  report ": WRAD1 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD0_delayed) = 'X') and (TO_X01(WRAD0_previous) /= 'X') then
		  assert false
		  report ": WRAD0 unknown"
		  severity Warning;
		end if;
	      else 
		RAM_TMP(WADDR) <= WD7_delayed & WD6_delayed & WD5_delayed & 
                                  WD4_delayed & WD3_delayed & WD2_delayed &
                                  WD1_delayed & WD0_delayed ; 
	      end if;
	    else
	      null;
	    end if;
	  when others =>
            if (TO_X01(WEN_previous) /= 'X') then
	      assert false
	      report ": WEN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      -- Convert Read Address Signal to Integer
      RADDR := ((INT(RDAD4_ipd)*16)+(INT(RDAD3_ipd)*8)+
		(INT(RDAD2_ipd)*4)+(INT(RDAD1_ipd)*2)+(INT(RDAD0_ipd)));

      if (RADDR < 0) then
	RD7_zd := 'X';
	RD6_zd := 'X';
	RD5_zd := 'X';
	RD4_zd := 'X';
	RD3_zd := 'X';
	RD2_zd := 'X';
	RD1_zd := 'X';
	RD0_zd := 'X';
	if (TO_X01(RDAD4_ipd) = 'X') and (TO_X01(RDAD4_previous) /= 'X') then
	  assert false
	  report ": RDAD4 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD3_ipd) = 'X') and (TO_X01(RDAD3_previous) /= 'X') then
	  assert false
	  report ": RDAD3 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD2_ipd) = 'X') and (TO_X01(RDAD2_previous) /= 'X') then
	  assert false
	  report ": RDAD2 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD1_ipd) = 'X') and (TO_X01(RDAD1_previous) /= 'X') then
	  assert false
	  report ": RDAD1 unknown"
	  severity Warning;
	end if;
	if (TO_X01(RDAD0_ipd) = 'X') and (TO_X01(RDAD0_previous) /= 'X') then
	  assert false
	  report ": RDAD0 unknown"
	  severity Warning;
	end if;
      else
	RD7_zd := RAM_TMP(RADDR)(7);
	RD6_zd := RAM_TMP(RADDR)(6);
	RD5_zd := RAM_TMP(RADDR)(5);
	RD4_zd := RAM_TMP(RADDR)(4);
	RD3_zd := RAM_TMP(RADDR)(3);
	RD2_zd := RAM_TMP(RADDR)(2);
	RD1_zd := RAM_TMP(RADDR)(1);
	RD0_zd := RAM_TMP(RADDR)(0);
      end if;
      
      WCLK_previous := WCLK_ipd;
      WEN_previous := WEN_delayed;
      WEN_delayed := WEN_ipd;
      BLKEN_previous := BLKEN_delayed;
      BLKEN_delayed := BLKEN_ipd;
      WD7_delayed := WD7_ipd;
      WD6_delayed := WD6_ipd;
      WD5_delayed := WD5_ipd;
      WD4_delayed := WD4_ipd;
      WD3_delayed := WD3_ipd;
      WD2_delayed := WD2_ipd;
      WD1_delayed := WD1_ipd;
      WD0_delayed := WD0_ipd;
      WRAD4_previous := WRAD4_delayed;
      WRAD3_previous := WRAD3_delayed;
      WRAD2_previous := WRAD2_delayed;
      WRAD1_previous := WRAD1_delayed;
      WRAD0_previous := WRAD0_delayed;
      WRAD4_delayed := WRAD4_ipd;
      WRAD3_delayed := WRAD3_ipd;
      WRAD2_delayed := WRAD2_ipd;
      WRAD1_delayed := WRAD1_ipd;
      WRAD0_delayed := WRAD0_ipd;
      RDAD4_previous := RDAD4_ipd;
      RDAD3_previous := RDAD3_ipd;
      RDAD2_previous := RDAD2_ipd;
      RDAD1_previous := RDAD1_ipd;
      RDAD0_previous := RDAD0_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD7,
	GlitchData => RD7_GlitchData,
	OutSignalName => "RD7",
	OutTemp => RD7_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD7), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD7), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD7), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD7), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD7), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD7), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD7), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD7), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD7), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD7), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD7), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD7), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD7), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD7), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD7), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD7), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD7), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD7), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD7), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD7), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD7), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD7), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD7), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD7), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD7), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD6,
	GlitchData => RD6_GlitchData,
	OutSignalName => "RD6",
	OutTemp => RD6_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD6), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD6), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD6), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD6), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD6), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD6), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD6), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD6), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD6), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD6), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD6), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD6), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD6), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD6), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD6), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD6), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD6), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD6), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD6), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD6), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD6), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD6), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD6), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD6), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD6), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD5,
	GlitchData => RD5_GlitchData,
	OutSignalName => "RD5",
	OutTemp => RD5_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD5), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD5), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD5), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD5), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD5), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD5), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD5), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD5), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD5), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD5), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD5), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD5), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD5), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD5), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD5), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD5), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD5), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD5), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD5), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD5), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD5), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD5), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD5), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD5), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD5), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD4,
	GlitchData => RD4_GlitchData,
	OutSignalName => "RD4",
	OutTemp => RD4_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD4), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD4), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD4), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD4), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD4), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD4), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD4), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD4), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD4), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD4), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD4), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD4), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD4), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD4), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD4), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD4), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD4), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD4), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD4), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD4), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD4), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD4), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD4), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD4), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD4), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD3,
	GlitchData => RD3_GlitchData,
	OutSignalName => "RD3",
	OutTemp => RD3_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD3), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD3), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD3), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD3), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD3), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD2,
	GlitchData => RD2_GlitchData,
	OutSignalName => "RD2",
	OutTemp => RD2_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD2), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD2), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD2), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD2), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD2), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD1,
	GlitchData => RD1_GlitchData,
	OutSignalName => "RD1",
	OutTemp => RD1_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD1), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD1), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD1), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD1), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD1), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD0,
	GlitchData => RD0_GlitchData,
	OutSignalName => "RD0",
	OutTemp => RD0_zd,
	Paths => (0 => (RDAD4_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
		  1 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
		  2 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
		  3 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
		  4 => (RDAD4_ipd'last_event,
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  5 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  6 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  7 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  8 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  9 => (RDAD3_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  10 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  11 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  12 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  13 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  14 => (RDAD2_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  15 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  16 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  17 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  18 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  19 => (RDAD1_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE),
                  20 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD4_RD0), TRUE),
                  21 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD3_RD0), TRUE),
                  22 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD2_RD0), TRUE),
                  23 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD1_RD0), TRUE),
                  24 => (RDAD0_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RDAD0_RD0), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

  end process VITALBehavior;

end VITAL_ACT;
-----------------------------------------------------------------
--  Proxy Modeling, Inc. 
--
--  Actel RAM8RF VHDL behavioral model
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - Jan/22/96 - Initial Delivery
-- 1.1 - 12/6/96 by DNW - Modified SL_TO_INT.
-- 1.2 - 3/3/97 by DNW - WDx_delayed variables added.
-- 1.3 - 3/6/98 by DNW - Issue "unknown" msg. only if 0/1->X Xtion.
-- 1.4 - 5/27/98 by DNW - Initaialize _ipd signals to X instead of 0.
-- 
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity RAM8RF is
  GENERIC (
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD7      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD6      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD5      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD4      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD4_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_negedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_negedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_negedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_negedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC;
        RD6    : OUT STD_ULOGIC;
        RD5    : OUT STD_ULOGIC;
        RD4    : OUT STD_ULOGIC;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of RAM8RF : entity is TRUE;
  
end RAM8RF;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM8RF is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal WRAD4_ipd : std_ulogic := 'X';
  signal WRAD3_ipd : std_ulogic := 'X';
  signal WRAD2_ipd : std_ulogic := 'X';
  signal WRAD1_ipd : std_ulogic := 'X';
  signal WRAD0_ipd : std_ulogic := 'X';
  signal WD7_ipd : std_ulogic := 'X';
  signal WD6_ipd : std_ulogic := 'X';
  signal WD5_ipd : std_ulogic := 'X';
  signal WD4_ipd : std_ulogic := 'X';
  signal WD3_ipd : std_ulogic := 'X';
  signal WD2_ipd : std_ulogic := 'X';
  signal WD1_ipd : std_ulogic := 'X';
  signal WD0_ipd : std_ulogic := 'X';
  signal RDAD4_ipd : std_ulogic := 'X';
  signal RDAD3_ipd : std_ulogic := 'X';
  signal RDAD2_ipd : std_ulogic := 'X';
  signal RDAD1_ipd : std_ulogic := 'X';
  signal RDAD0_ipd : std_ulogic := 'X';
  signal BLKEN_ipd : std_ulogic := 'X';
  signal WEN_ipd : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal REN_ipd : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  type MEM is array(0 to 31) of std_ulogic_vector(7 downto 0);
   signal RAM_TMP : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (WRAD4_ipd, WRAD4, VitalExtendToFillDelay(tipd_WRAD4));
    VitalWireDelay (WRAD3_ipd, WRAD3, VitalExtendToFillDelay(tipd_WRAD3));
    VitalWireDelay (WRAD2_ipd, WRAD2, VitalExtendToFillDelay(tipd_WRAD2));
    VitalWireDelay (WRAD1_ipd, WRAD1, VitalExtendToFillDelay(tipd_WRAD1));
    VitalWireDelay (WRAD0_ipd, WRAD0, VitalExtendToFillDelay(tipd_WRAD0));
    VitalWireDelay (WD7_ipd, WD7, VitalExtendToFillDelay(tipd_WD7));
    VitalWireDelay (WD6_ipd, WD6, VitalExtendToFillDelay(tipd_WD6));
    VitalWireDelay (WD5_ipd, WD5, VitalExtendToFillDelay(tipd_WD5));
    VitalWireDelay (WD4_ipd, WD4, VitalExtendToFillDelay(tipd_WD4));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (RDAD4_ipd, RDAD4, VitalExtendToFillDelay(tipd_RDAD4));
    VitalWireDelay (RDAD3_ipd, RDAD3, VitalExtendToFillDelay(tipd_RDAD3));
    VitalWireDelay (RDAD2_ipd, RDAD2, VitalExtendToFillDelay(tipd_RDAD2));
    VitalWireDelay (RDAD1_ipd, RDAD1, VitalExtendToFillDelay(tipd_RDAD1));
    VitalWireDelay (RDAD0_ipd, RDAD0, VitalExtendToFillDelay(tipd_RDAD0));
    VitalWireDelay (BLKEN_ipd, BLKEN, VitalExtendToFillDelay(tipd_BLKEN));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (REN_ipd, REN, VitalExtendToFillDelay(tipd_REN));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (RDAD4_ipd, RDAD3_ipd, RDAD2_ipd, RDAD1_ipd, 
		RDAD0_ipd, REN_ipd, RCLK_ipd, WD7_ipd, WD6_ipd, WD5_ipd, 
		WD4_ipd, WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd, WRAD4_ipd, 
		WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, WEN_ipd, 
		BLKEN_ipd, BLKENS, WCLK_ipd)

     --  Read Timing Check Results
     variable Tviol_RDAD4_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD4_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD3_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD3_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD2_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD2_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD1_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD1_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD0_RCLK_negedge : X01 := '0';
     variable TmDt_RDAD0_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_REN_RCLK_negedge : X01 := '0';
     variable TmDt_REN_RCLK_negedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_WD7_WCLK_posedge : X01 := '0';
     variable TmDt_WD7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD6_WCLK_posedge : X01 := '0';
     variable TmDt_WD6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD5_WCLK_posedge : X01 := '0';
     variable TmDt_WD5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD4_WCLK_posedge : X01 := '0';
     variable TmDt_WD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD3_WCLK_posedge : X01 := '0';
     variable TmDt_WD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_posedge : X01 := '0';
     variable TmDt_WD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_posedge : X01 := '0';
     variable TmDt_WD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_posedge : X01 := '0';
     variable TmDt_WD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD4_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD3_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD2_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD1_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD0_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_posedge : X01 := '0';
     variable TmDt_WEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_BLKEN_WCLK_posedge : X01 := '0';
     variable TmDt_BLKEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     --type SL_TO_INT is array(std_ulogic range <>) of integer;
     --constant INT :SL_TO_INT('U' to '-') := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     variable RD7_zd : std_ulogic;
     variable RD6_zd : std_ulogic;
     variable RD5_zd : std_ulogic;
     variable RD4_zd : std_ulogic;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD7_GlitchData : VitalGlitchDataType;
     variable RD6_GlitchData : VitalGlitchDataType;
     variable RD5_GlitchData : VitalGlitchDataType;
     variable RD4_GlitchData : VitalGlitchDataType;
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;
  
     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable WEN_delayed : std_ulogic := 'X';
     variable REN_delayed : std_ulogic := 'X';
     variable WEN_previous : std_ulogic := 'X';
     variable REN_previous : std_ulogic := 'X';
     variable BLKEN_delayed : std_ulogic := 'X';
     variable BLKEN_previous : std_ulogic := 'X';
     variable WD7_delayed : std_ulogic := 'X';
     variable WD6_delayed : std_ulogic := 'X';
     variable WD5_delayed : std_ulogic := 'X';
     variable WD4_delayed : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WRAD4_delayed : std_ulogic := 'X';
     variable WRAD3_delayed : std_ulogic := 'X';
     variable WRAD2_delayed : std_ulogic := 'X';
     variable WRAD1_delayed : std_ulogic := 'X';
     variable WRAD0_delayed : std_ulogic := 'X';
     variable WRAD4_previous : std_ulogic := 'X';
     variable WRAD3_previous : std_ulogic := 'X';
     variable WRAD2_previous : std_ulogic := 'X';
     variable WRAD1_previous : std_ulogic := 'X';
     variable WRAD0_previous : std_ulogic := 'X';
     variable RDAD4_delayed : std_ulogic := 'X';
     variable RDAD3_delayed : std_ulogic := 'X';
     variable RDAD2_delayed : std_ulogic := 'X';
     variable RDAD1_delayed : std_ulogic := 'X';
     variable RDAD0_delayed : std_ulogic := 'X';
     variable RDAD4_previous : std_ulogic := 'X';
     variable RDAD3_previous : std_ulogic := 'X';
     variable RDAD2_previous : std_ulogic := 'X';
     variable RDAD1_previous : std_ulogic := 'X';
     variable RDAD0_previous : std_ulogic := 'X';
  
  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RDAD high or low before RCLK falling
      --   Hold  RDAD high or low after RCLK falling

      VitalSetupHoldCheck ( Tviol_RDAD4_RCLK_negedge,
                            TmDt_RDAD4_RCLK_negedge,
                            RDAD4_ipd, "RDAD4",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD4_RCLK_noedge_negedge,
                            tsetup_RDAD4_RCLK_noedge_negedge,
                            thold_RDAD4_RCLK_noedge_negedge,
                            thold_RDAD4_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD3_RCLK_negedge,
                            TmDt_RDAD3_RCLK_negedge,
                            RDAD3_ipd, "RDAD3",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD3_RCLK_noedge_negedge,
                            tsetup_RDAD3_RCLK_noedge_negedge,
                            thold_RDAD3_RCLK_noedge_negedge,
                            thold_RDAD3_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD2_RCLK_negedge,
                            TmDt_RDAD2_RCLK_negedge,
                            RDAD2_ipd, "RDAD2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD2_RCLK_noedge_negedge,
                            tsetup_RDAD2_RCLK_noedge_negedge,
                            thold_RDAD2_RCLK_noedge_negedge,
                            thold_RDAD2_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD1_RCLK_negedge,
                            TmDt_RDAD1_RCLK_negedge,
                            RDAD1_ipd, "RDAD1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD1_RCLK_noedge_negedge,
                            tsetup_RDAD1_RCLK_noedge_negedge,
                            thold_RDAD1_RCLK_noedge_negedge,
                            thold_RDAD1_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD0_RCLK_negedge,
                            TmDt_RDAD0_RCLK_negedge,
                            RDAD0_ipd, "RDAD0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD0_RCLK_noedge_negedge,
                            tsetup_RDAD0_RCLK_noedge_negedge,
                            thold_RDAD0_RCLK_noedge_negedge,
                            thold_RDAD0_RCLK_noedge_negedge,
                            (To_X01(REN_ipd)='1'),
                            '\',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup REN high before RCLK falling
      --   Hold  REN high after RCLK falling

      VitalSetupHoldCheck ( Tviol_REN_RCLK_negedge,
                            TmDt_REN_RCLK_negedge,
                            REN_ipd, "REN",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_REN_RCLK_noedge_negedge,
                            tsetup_REN_RCLK_noedge_negedge,
                            thold_REN_RCLK_noedge_negedge,
                            thold_REN_RCLK_noedge_negedge,
                            TimingCheckOn,
                            '\',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup BLKEN high or low before WCLK rising
      --   Hold  BLKEN high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_BLKEN_WCLK_posedge,
                            TmDt_BLKEN_WCLK_posedge,
                            BLKEN_ipd, "BLKEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_BLKEN_WCLK_noedge_posedge,
                            tsetup_BLKEN_WCLK_noedge_posedge,
                            thold_BLKEN_WCLK_noedge_posedge,
                            thold_BLKEN_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WRAD high or low before WCLK rising
      --   Hold  WRAD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WRAD4_WCLK_posedge,
                            TmDt_WRAD4_WCLK_posedge,
                            WRAD4_ipd, "WRAD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD4_WCLK_noedge_posedge,
                            tsetup_WRAD4_WCLK_noedge_posedge,
                            thold_WRAD4_WCLK_noedge_posedge,
                            thold_WRAD4_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD3_WCLK_posedge,
                            TmDt_WRAD3_WCLK_posedge,
                            WRAD3_ipd, "WRAD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD3_WCLK_noedge_posedge,
                            tsetup_WRAD3_WCLK_noedge_posedge,
                            thold_WRAD3_WCLK_noedge_posedge,
                            thold_WRAD3_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD2_WCLK_posedge,
                            TmDt_WRAD2_WCLK_posedge,
                            WRAD2_ipd, "WRAD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD2_WCLK_noedge_posedge,
                            tsetup_WRAD2_WCLK_noedge_posedge,
                            thold_WRAD2_WCLK_noedge_posedge,
                            thold_WRAD2_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD1_WCLK_posedge,
                            TmDt_WRAD1_WCLK_posedge,
                            WRAD1_ipd, "WRAD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD1_WCLK_noedge_posedge,
                            tsetup_WRAD1_WCLK_noedge_posedge,
                            thold_WRAD1_WCLK_noedge_posedge,
                            thold_WRAD1_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD0_WCLK_posedge,
                            TmDt_WRAD0_WCLK_posedge,
                            WRAD0_ipd, "WRAD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD0_WCLK_noedge_posedge,
                            tsetup_WRAD0_WCLK_noedge_posedge,
                            thold_WRAD0_WCLK_noedge_posedge,
                            thold_WRAD0_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WD high or low before WCLK rising
      --   Hold  WD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WD7_WCLK_posedge,
                            TmDt_WD7_WCLK_posedge,
                            WD7_ipd, "WD7",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD7_WCLK_noedge_posedge,
                            tsetup_WD7_WCLK_noedge_posedge,
                            thold_WD7_WCLK_noedge_posedge,
                            thold_WD7_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD6_WCLK_posedge,
                            TmDt_WD6_WCLK_posedge,
                            WD6_ipd, "WD6",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD6_WCLK_noedge_posedge,
                            tsetup_WD6_WCLK_noedge_posedge,
                            thold_WD6_WCLK_noedge_posedge,
                            thold_WD6_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD5_WCLK_posedge,
                            TmDt_WD5_WCLK_posedge,
                            WD5_ipd, "WD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD5_WCLK_noedge_posedge,
                            tsetup_WD5_WCLK_noedge_posedge,
                            thold_WD5_WCLK_noedge_posedge,
                            thold_WD5_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD4_WCLK_posedge,
                            TmDt_WD4_WCLK_posedge,
                            WD4_ipd, "WD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD4_WCLK_noedge_posedge,
                            tsetup_WD4_WCLK_noedge_posedge,
                            thold_WD4_WCLK_noedge_posedge,
                            thold_WD4_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_posedge,
                            TmDt_WD3_WCLK_posedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_noedge_posedge,
                            tsetup_WD3_WCLK_noedge_posedge,
                            thold_WD3_WCLK_noedge_posedge,
                            thold_WD3_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_posedge,
                            TmDt_WD2_WCLK_posedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_noedge_posedge,
                            tsetup_WD2_WCLK_noedge_posedge,
                            thold_WD2_WCLK_noedge_posedge,
                            thold_WD2_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_posedge,
                            TmDt_WD1_WCLK_posedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_noedge_posedge,
                            tsetup_WD1_WCLK_noedge_posedge,
                            thold_WD1_WCLK_noedge_posedge,
                            thold_WD1_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_posedge,
                            TmDt_WD0_WCLK_posedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_noedge_posedge,
                            tsetup_WD0_WCLK_noedge_posedge,
                            thold_WD0_WCLK_noedge_posedge,
                            thold_WD0_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup WEN high before WCLK rising
      --   Hold  WEN high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_posedge,
                            TmDt_WEN_WCLK_posedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_noedge_posedge,
                            tsetup_WEN_WCLK_noedge_posedge,
                            thold_WEN_WCLK_noedge_posedge,
                            thold_WEN_WCLK_noedge_posedge,
                            (To_X01(BLKEN_ipd)=BLKENS),
                            '/',
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM8RF",
                            TRUE,
                            TRUE,
                            ERROR
                            );
    
    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      -- Convert Write Address Signal to Integer
      WADDR := ((INT(WRAD4_delayed)*16)+(INT(WRAD3_delayed)*8)+(INT(WRAD2_delayed)*4)
		+(INT(WRAD1_delayed)*2)+(INT(WRAD0_delayed)));

      if (TO_X01(WCLK_ipd)='X') then
        if (TO_X01(WCLK_previous) /= 'X') then
	  assert false
	  report ": WCLK unknown"
	  severity Warning;
	end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	case TO_X01(WEN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (TO_X01(BLKEN_delayed) = 'X') then
              if (TO_X01(BLKEN_previous) /= 'X') then
	        assert false
	        report ": BLKEN unknown"
	        severity Warning;
	      end if;
	    elsif (TO_X01(BLKEN_delayed) = BLKENS) then
	      if (WADDR < 0) then
		if (TO_X01(WRAD4_delayed) = 'X') and (TO_X01(WRAD4_previous) /= 'X') then
		  assert false
		  report ": WRAD4 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD3_delayed) = 'X') and (TO_X01(WRAD3_previous) /= 'X') then
		  assert false
		  report ": WRAD3 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD2_delayed) = 'X') and (TO_X01(WRAD2_previous) /= 'X') then
		  assert false
		  report ": WRAD2 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD1_delayed) = 'X') and (TO_X01(WRAD1_previous) /= 'X') then
		  assert false
		  report ": WRAD1 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD0_delayed) = 'X') and (TO_X01(WRAD0_previous) /= 'X') then
		  assert false
		  report ": WRAD0 unknown"
		  severity Warning;
		end if;
	      else 
		RAM_TMP(WADDR) <= WD7_delayed & WD6_delayed & WD5_delayed & 
                                  WD4_delayed & WD3_delayed & WD2_delayed &
                                  WD1_delayed & WD0_delayed ; 
	      end if;
	    else
	      null;
	    end if;
	  when others =>
            if (TO_X01(WEN_previous) /= 'X') then
	      assert false
	      report ": WEN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      -- Convert Read Address Signal to Integer
      RADDR := ((INT(RDAD4_delayed)*16)+(INT(RDAD3_delayed)*8)+(INT(RDAD2_delayed)*4)
		+(INT(RDAD1_delayed)*2)+(INT(RDAD0_delayed)));

      if (TO_X01(RCLK_ipd) = 'X') then
	RD7_zd := 'X';
	RD6_zd := 'X';
	RD5_zd := 'X';
	RD4_zd := 'X';
	RD3_zd := 'X';
	RD2_zd := 'X';
	RD1_zd := 'X';
	RD0_zd := 'X';
	if (TO_X01(RCLK_previous) /= 'X') then
	  assert false
	  report ": RCLK unknown"
	  severity Warning;
	end if;
      elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '0')) then
	case TO_X01(REN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (RADDR < 0) then
	      RD7_zd := 'X';
	      RD6_zd := 'X';
	      RD5_zd := 'X';
	      RD4_zd := 'X';
	      RD3_zd := 'X';
	      RD2_zd := 'X';
	      RD1_zd := 'X';
	      RD0_zd := 'X';
	      if (TO_X01(RDAD4_delayed) = 'X') and (TO_X01(RDAD4_previous) /= 'X') then
		assert false
		report ": RDAD4 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD3_delayed) = 'X') and (TO_X01(RDAD3_previous) /= 'X') then
		assert false
		report ": RDAD3 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD2_delayed) = 'X') and (TO_X01(RDAD2_previous) /= 'X') then
		assert false
		report ": RDAD2 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD1_delayed) = 'X') and (TO_X01(RDAD1_previous) /= 'X') then
		assert false
		report ": RDAD1 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD0_delayed) = 'X') and (TO_X01(RDAD0_previous) /= 'X') then
		assert false
		report ": RDAD0 unknown"
		severity Warning;
	      end if;
	    else
	      RD7_zd := RAM_TMP(RADDR)(7);
	      RD6_zd := RAM_TMP(RADDR)(6);
	      RD5_zd := RAM_TMP(RADDR)(5);
	      RD4_zd := RAM_TMP(RADDR)(4);
	      RD3_zd := RAM_TMP(RADDR)(3);
	      RD2_zd := RAM_TMP(RADDR)(2);
	      RD1_zd := RAM_TMP(RADDR)(1);
	      RD0_zd := RAM_TMP(RADDR)(0);
	    end if;
	  when others =>
	    RD7_zd := 'X';
	    RD6_zd := 'X';
	    RD5_zd := 'X';
	    RD4_zd := 'X';
	    RD3_zd := 'X';
	    RD2_zd := 'X';
	    RD1_zd := 'X';
	    RD0_zd := 'X';
            if (TO_X01(REN_previous) /= 'X') then
	      assert false
	      report ": REN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;
      
      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      WEN_previous := WEN_delayed;
      REN_previous := REN_delayed;
      WEN_delayed := WEN_ipd;
      REN_delayed := REN_ipd;
      BLKEN_previous := BLKEN_delayed;
      BLKEN_delayed := BLKEN_ipd;
      WD7_delayed := WD7_ipd;
      WD6_delayed := WD6_ipd;
      WD5_delayed := WD5_ipd;
      WD4_delayed := WD4_ipd;
      WD3_delayed := WD3_ipd;
      WD2_delayed := WD2_ipd;
      WD1_delayed := WD1_ipd;
      WD0_delayed := WD0_ipd;
      WRAD4_previous := WRAD4_delayed;
      WRAD3_previous := WRAD3_delayed;
      WRAD2_previous := WRAD2_delayed;
      WRAD1_previous := WRAD1_delayed;
      WRAD0_previous := WRAD0_delayed;
      WRAD4_delayed := WRAD4_ipd;
      WRAD3_delayed := WRAD3_ipd;
      WRAD2_delayed := WRAD2_ipd;
      WRAD1_delayed := WRAD1_ipd;
      WRAD0_delayed := WRAD0_ipd;
      RDAD4_previous := RDAD4_delayed;
      RDAD3_previous := RDAD3_delayed;
      RDAD2_previous := RDAD2_delayed;
      RDAD1_previous := RDAD1_delayed;
      RDAD0_previous := RDAD0_delayed;
      RDAD4_delayed := RDAD4_ipd;
      RDAD3_delayed := RDAD3_ipd;
      RDAD2_delayed := RDAD2_ipd;
      RDAD1_delayed := RDAD1_ipd;
      RDAD0_delayed := RDAD0_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD7,
	GlitchData => RD7_GlitchData,
	OutSignalName => "RD7",
	OutTemp => RD7_zd,
	Paths => (0 => (RCLK_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RCLK_RD7), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD6,
	GlitchData => RD6_GlitchData,
	OutSignalName => "RD6",
	OutTemp => RD6_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD6), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD5,
	GlitchData => RD5_GlitchData,
	OutSignalName => "RD5",
	OutTemp => RD5_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD5), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD4,
	GlitchData => RD4_GlitchData,
	OutSignalName => "RD4",
	OutTemp => RD4_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD4), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD3,
	GlitchData => RD3_GlitchData,
	OutSignalName => "RD3",
	OutTemp => RD3_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD3), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD2,
	GlitchData => RD2_GlitchData,
	OutSignalName => "RD2",
	OutTemp => RD2_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD2), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD1,
	GlitchData => RD1_GlitchData,
	OutSignalName => "RD1",
	OutTemp => RD1_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD1), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD0,
	GlitchData => RD0_GlitchData,
	OutSignalName => "RD0",
	OutTemp => RD0_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD0), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

  end process VITALBehavior;

end VITAL_ACT;
-----------------------------------------------------------------
--  Proxy Modeling, Inc. 
--
--  Actel RAM8RR VHDL behavioral model
--  Uses VITAL95 package
--
-- =================
-- Revision History
-- =================
--
-- 1.0 - Jan/22/96 - Initial Delivery
-- 1.1 - 12/6/96 by DNW - Modified SL_TO_INT.
-- 1.2 - 3/3/97 by DNW - WDx_delayed variables added.
-- 1.3 - 3/6/98 by DNW - Issue "unknown" msg. only if 0/1->X Xtion.
-- 1.4 - 5/27/98 by DNW - Initaialize _ipd signals to X instead of 0.
-- 
-----------------------------------------------------------------

LIBRARY IEEE;
  use IEEE.STD_LOGIC_1164.all;
  use IEEE.VITAL_timing.all;

-- #########################################################
-- # ENTITY declaration
-- #########################################################
  
entity RAM8RR is
  GENERIC (
        tipd_RDAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RDAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_REN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_RCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD7      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD6      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD5      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD4      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD3      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD2      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD1      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WD0      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD4    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD3    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD2    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD1    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WRAD0    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WEN      : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_BLKEN    : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tipd_WCLK     : VitalDelayType01 := (1.000 ns, 1.000 ns);
        tpd_RCLK_RD7 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD6 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD5 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD4 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD3 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD2 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD1 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tpd_RCLK_RD0 : VitalDelayType01 := (0.000 ns, 0.000 ns);
        tsetup_RDAD4_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD3_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD2_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD1_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_RDAD0_RCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD4_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD3_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD2_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD1_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WRAD0_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tsetup_WD7_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD6_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD5_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD4_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD3_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD2_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD1_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WD0_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        thold_RDAD4_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD3_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD2_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD1_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_RDAD0_RCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD4_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD3_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD2_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD1_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WRAD0_WCLK_noedge_posedge    : VitalDelayType := 0.000 ns;
        thold_WD7_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD6_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD5_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD4_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD3_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD2_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD1_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WD0_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        tsetup_REN_RCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
        tsetup_WEN_WCLK_noedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        thold_REN_RCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
        thold_WEN_WCLK_noedge_posedge      : VitalDelayType := 0.000 ns;
	thold_BLKEN_WCLK_noedge_posedge   : VitalDelayType := 0.000 ns;
        tpw_RCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_RCLK_negedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_posedge    : VitalDelayType := 0.000 ns;
        tpw_WCLK_negedge    : VitalDelayType := 0.000 ns;
        TimingCheckOn : BOOLEAN := TRUE;
        InstancePath  : STRING := "*"
        );
  PORT (
        WRAD4  : IN STD_ULOGIC ;
        WRAD3  : IN STD_ULOGIC ;
        WRAD2  : IN STD_ULOGIC ;
        WRAD1  : IN STD_ULOGIC ;
        WRAD0  : IN STD_ULOGIC ;
        WD7    : IN STD_ULOGIC ;
        WD6    : IN STD_ULOGIC ;
        WD5    : IN STD_ULOGIC ;
        WD4    : IN STD_ULOGIC ;
        WD3    : IN STD_ULOGIC ;
        WD2    : IN STD_ULOGIC ;
        WD1    : IN STD_ULOGIC ;
        WD0    : IN STD_ULOGIC ;
        RDAD4  : IN STD_ULOGIC ;
        RDAD3  : IN STD_ULOGIC ;
        RDAD2  : IN STD_ULOGIC ;
        RDAD1  : IN STD_ULOGIC ;
        RDAD0  : IN STD_ULOGIC ;
        BLKEN  : IN STD_ULOGIC ;
        BLKENS : IN STD_ULOGIC ;
        WEN    : IN STD_ULOGIC ;
        WCLK   : IN STD_ULOGIC ;
        REN    : IN STD_ULOGIC ;
        RCLK   : IN STD_ULOGIC ;
        RD7    : OUT STD_ULOGIC;
        RD6    : OUT STD_ULOGIC;
        RD5    : OUT STD_ULOGIC;
        RD4    : OUT STD_ULOGIC;
        RD3    : OUT STD_ULOGIC;
        RD2    : OUT STD_ULOGIC;
        RD1    : OUT STD_ULOGIC;
        RD0    : OUT STD_ULOGIC
        );

  attribute VITAL_LEVEL0 of RAM8RR : entity is TRUE;
  
end RAM8RR;

-- #########################################################
-- # ARCHITECTURE declaration
-- #########################################################
architecture VITAL_ACT of RAM8RR is

  attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

  signal WRAD4_ipd : std_ulogic := 'X';
  signal WRAD3_ipd : std_ulogic := 'X';
  signal WRAD2_ipd : std_ulogic := 'X';
  signal WRAD1_ipd : std_ulogic := 'X';
  signal WRAD0_ipd : std_ulogic := 'X';
  signal WD7_ipd : std_ulogic := 'X';
  signal WD6_ipd : std_ulogic := 'X';
  signal WD5_ipd : std_ulogic := 'X';
  signal WD4_ipd : std_ulogic := 'X';
  signal WD3_ipd : std_ulogic := 'X';
  signal WD2_ipd : std_ulogic := 'X';
  signal WD1_ipd : std_ulogic := 'X';
  signal WD0_ipd : std_ulogic := 'X';
  signal RDAD4_ipd : std_ulogic := 'X';
  signal RDAD3_ipd : std_ulogic := 'X';
  signal RDAD2_ipd : std_ulogic := 'X';
  signal RDAD1_ipd : std_ulogic := 'X';
  signal RDAD0_ipd : std_ulogic := 'X';
  signal BLKEN_ipd : std_ulogic := 'X';
  signal WEN_ipd : std_ulogic := 'X';
  signal WCLK_ipd : std_ulogic := 'X';
  signal REN_ipd : std_ulogic := 'X';
  signal RCLK_ipd : std_ulogic := 'X';
  type MEM is array(0 to 31) of std_ulogic_vector(7 downto 0);
   signal RAM_TMP : MEM;
  
begin  --  VITAL_ACT 

  -- #########################################################
  -- # INPUT PATH DELAYS
  -- #########################################################

  WIRE_DELAY: block
  
  begin  --  block WIRE_DELAY 
    VitalWireDelay (WRAD4_ipd, WRAD4, VitalExtendToFillDelay(tipd_WRAD4));
    VitalWireDelay (WRAD3_ipd, WRAD3, VitalExtendToFillDelay(tipd_WRAD3));
    VitalWireDelay (WRAD2_ipd, WRAD2, VitalExtendToFillDelay(tipd_WRAD2));
    VitalWireDelay (WRAD1_ipd, WRAD1, VitalExtendToFillDelay(tipd_WRAD1));
    VitalWireDelay (WRAD0_ipd, WRAD0, VitalExtendToFillDelay(tipd_WRAD0));
    VitalWireDelay (WD7_ipd, WD7, VitalExtendToFillDelay(tipd_WD7));
    VitalWireDelay (WD6_ipd, WD6, VitalExtendToFillDelay(tipd_WD6));
    VitalWireDelay (WD5_ipd, WD5, VitalExtendToFillDelay(tipd_WD5));
    VitalWireDelay (WD4_ipd, WD4, VitalExtendToFillDelay(tipd_WD4));
    VitalWireDelay (WD3_ipd, WD3, VitalExtendToFillDelay(tipd_WD3));
    VitalWireDelay (WD2_ipd, WD2, VitalExtendToFillDelay(tipd_WD2));
    VitalWireDelay (WD1_ipd, WD1, VitalExtendToFillDelay(tipd_WD1));
    VitalWireDelay (WD0_ipd, WD0, VitalExtendToFillDelay(tipd_WD0));
    VitalWireDelay (RDAD4_ipd, RDAD4, VitalExtendToFillDelay(tipd_RDAD4));
    VitalWireDelay (RDAD3_ipd, RDAD3, VitalExtendToFillDelay(tipd_RDAD3));
    VitalWireDelay (RDAD2_ipd, RDAD2, VitalExtendToFillDelay(tipd_RDAD2));
    VitalWireDelay (RDAD1_ipd, RDAD1, VitalExtendToFillDelay(tipd_RDAD1));
    VitalWireDelay (RDAD0_ipd, RDAD0, VitalExtendToFillDelay(tipd_RDAD0));
    VitalWireDelay (BLKEN_ipd, BLKEN, VitalExtendToFillDelay(tipd_BLKEN));
    VitalWireDelay (WEN_ipd, WEN, VitalExtendToFillDelay(tipd_WEN));
    VitalWireDelay (WCLK_ipd, WCLK, VitalExtendToFillDelay(tipd_WCLK));
    VitalWireDelay (REN_ipd, REN, VitalExtendToFillDelay(tipd_REN));
    VitalWireDelay (RCLK_ipd, RCLK, VitalExtendToFillDelay(tipd_RCLK));
  end block WIRE_DELAY;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  VITALBehavior : process (RDAD4_ipd, RDAD3_ipd, RDAD2_ipd, RDAD1_ipd, 
		RDAD0_ipd, REN_ipd, RCLK_ipd, WD7_ipd, WD6_ipd, WD5_ipd, 
		WD4_ipd, WD3_ipd, WD2_ipd, WD1_ipd, WD0_ipd, WRAD4_ipd, 
		WRAD3_ipd, WRAD2_ipd, WRAD1_ipd, WRAD0_ipd, WEN_ipd, 
		BLKEN_ipd, BLKENS, WCLK_ipd)

     --  Read Timing Check Results
     variable Tviol_RDAD4_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD4_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD3_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD3_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD2_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD2_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD1_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD1_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDAD0_RCLK_posedge : X01 := '0';
     variable TmDt_RDAD0_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_REN_RCLK_posedge : X01 := '0';
     variable TmDt_REN_RCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_RCLK : X01 := '0';
     variable PeriodData_RCLK : VitalPeriodDataType := VitalPeriodDataInit;
      
     --  Write Timing Check Results
     variable Tviol_WD7_WCLK_posedge : X01 := '0';
     variable TmDt_WD7_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD6_WCLK_posedge : X01 := '0';
     variable TmDt_WD6_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD5_WCLK_posedge : X01 := '0';
     variable TmDt_WD5_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD4_WCLK_posedge : X01 := '0';
     variable TmDt_WD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD3_WCLK_posedge : X01 := '0';
     variable TmDt_WD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD2_WCLK_posedge : X01 := '0';
     variable TmDt_WD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD1_WCLK_posedge : X01 := '0';
     variable TmDt_WD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WD0_WCLK_posedge : X01 := '0';
     variable TmDt_WD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD4_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD4_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD3_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD3_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD2_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD2_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD1_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD1_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRAD0_WCLK_posedge : X01 := '0';
     variable TmDt_WRAD0_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WEN_WCLK_posedge : X01 := '0';
     variable TmDt_WEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_BLKEN_WCLK_posedge : X01 := '0';
     variable TmDt_BLKEN_WCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
     variable Pviol_WCLK : X01 := '0';
     variable PeriodData_WCLK : VitalPeriodDataType := VitalPeriodDataInit;
                
     --  Functional Results
     --type SL_TO_INT is array(std_ulogic range <>) of integer;
     --constant INT :SL_TO_INT('U' to '-') := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);
     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     variable RD7_zd : std_ulogic;
     variable RD6_zd : std_ulogic;
     variable RD5_zd : std_ulogic;
     variable RD4_zd : std_ulogic;
     variable RD3_zd : std_ulogic;
     variable RD2_zd : std_ulogic;
     variable RD1_zd : std_ulogic;
     variable RD0_zd : std_ulogic;
      
     -- Output Glitch Detection Support Variables
     variable RD7_GlitchData : VitalGlitchDataType;
     variable RD6_GlitchData : VitalGlitchDataType;
     variable RD5_GlitchData : VitalGlitchDataType;
     variable RD4_GlitchData : VitalGlitchDataType;
     variable RD3_GlitchData : VitalGlitchDataType;
     variable RD2_GlitchData : VitalGlitchDataType;
     variable RD1_GlitchData : VitalGlitchDataType;
     variable RD0_GlitchData : VitalGlitchDataType;
  
     -- Last value variables
     variable WCLK_previous : std_ulogic := 'X';
     variable RCLK_previous : std_ulogic := 'X';
     variable WEN_delayed : std_ulogic := 'X';
     variable REN_delayed : std_ulogic := 'X';
     variable WEN_previous : std_ulogic := 'X';
     variable REN_previous : std_ulogic := 'X';
     variable BLKEN_delayed : std_ulogic := 'X';
     variable BLKEN_previous : std_ulogic := 'X';
     variable WD7_delayed : std_ulogic := 'X';
     variable WD6_delayed : std_ulogic := 'X';
     variable WD5_delayed : std_ulogic := 'X';
     variable WD4_delayed : std_ulogic := 'X';
     variable WD3_delayed : std_ulogic := 'X';
     variable WD2_delayed : std_ulogic := 'X';
     variable WD1_delayed : std_ulogic := 'X';
     variable WD0_delayed : std_ulogic := 'X';
     variable WRAD4_delayed : std_ulogic := 'X';
     variable WRAD3_delayed : std_ulogic := 'X';
     variable WRAD2_delayed : std_ulogic := 'X';
     variable WRAD1_delayed : std_ulogic := 'X';
     variable WRAD0_delayed : std_ulogic := 'X';
     variable WRAD4_previous : std_ulogic := 'X';
     variable WRAD3_previous : std_ulogic := 'X';
     variable WRAD2_previous : std_ulogic := 'X';
     variable WRAD1_previous : std_ulogic := 'X';
     variable WRAD0_previous : std_ulogic := 'X';
     variable RDAD4_delayed : std_ulogic := 'X';
     variable RDAD3_delayed : std_ulogic := 'X';
     variable RDAD2_delayed : std_ulogic := 'X';
     variable RDAD1_delayed : std_ulogic := 'X';
     variable RDAD0_delayed : std_ulogic := 'X';
     variable RDAD4_previous : std_ulogic := 'X';
     variable RDAD3_previous : std_ulogic := 'X';
     variable RDAD2_previous : std_ulogic := 'X';
     variable RDAD1_previous : std_ulogic := 'X';
     variable RDAD0_previous : std_ulogic := 'X';
  
  begin  --  process VITALBehavior 

    if (TimingCheckOn) then
      -- #########################################################
      -- # Read Timing Check Section
      -- #########################################################
    
      --   Setup RDAD high or low before RCLK rising
      --   Hold  RDAD high or low after RCLK rising

      VitalSetupHoldCheck ( Tviol_RDAD4_RCLK_posedge,
                            TmDt_RDAD4_RCLK_posedge,
                            RDAD4_ipd, "RDAD4",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD4_RCLK_noedge_posedge,
                            tsetup_RDAD4_RCLK_noedge_posedge,
                            thold_RDAD4_RCLK_noedge_posedge,
                            thold_RDAD4_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD3_RCLK_posedge,
                            TmDt_RDAD3_RCLK_posedge,
                            RDAD3_ipd, "RDAD3",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD3_RCLK_noedge_posedge,
                            tsetup_RDAD3_RCLK_noedge_posedge,
                            thold_RDAD3_RCLK_noedge_posedge,
                            thold_RDAD3_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD2_RCLK_posedge,
                            TmDt_RDAD2_RCLK_posedge,
                            RDAD2_ipd, "RDAD2",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD2_RCLK_noedge_posedge,
                            tsetup_RDAD2_RCLK_noedge_posedge,
                            thold_RDAD2_RCLK_noedge_posedge,
                            thold_RDAD2_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD1_RCLK_posedge,
                            TmDt_RDAD1_RCLK_posedge,
                            RDAD1_ipd, "RDAD1",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD1_RCLK_noedge_posedge,
                            tsetup_RDAD1_RCLK_noedge_posedge,
                            thold_RDAD1_RCLK_noedge_posedge,
                            thold_RDAD1_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_RDAD0_RCLK_posedge,
                            TmDt_RDAD0_RCLK_posedge,
                            RDAD0_ipd, "RDAD0",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_RDAD0_RCLK_noedge_posedge,
                            tsetup_RDAD0_RCLK_noedge_posedge,
                            thold_RDAD0_RCLK_noedge_posedge,
                            thold_RDAD0_RCLK_noedge_posedge,
                            (To_X01(REN_ipd)='1'),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup REN high before RCLK rising
      --   Hold  REN high after RCLK rising

      VitalSetupHoldCheck ( Tviol_REN_RCLK_posedge,
                            TmDt_REN_RCLK_posedge,
                            REN_ipd, "REN",
                            0.0 ns,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
                            tsetup_REN_RCLK_noedge_posedge,
			    tsetup_REN_RCLK_noedge_posedge,
                            thold_REN_RCLK_noedge_posedge,
                            thold_REN_RCLK_noedge_posedge,
                            TimingCheckOn,
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of RCLK 

      VitalPeriodPulseCheck ( Pviol_RCLK,
                            PeriodData_RCLK,
                            RCLK_ipd, "RCLK",
                            0.0 ns,
			    tpw_RCLK_posedge + tpw_RCLK_negedge,
                            tpw_RCLK_posedge,
                            tpw_RCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      -- #########################################################
      -- # Write Timing Check Section
      -- #########################################################

      --   Setup BLKEN high or low before WCLK rising
      --   Hold  BLKEN high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_BLKEN_WCLK_posedge,
                            TmDt_BLKEN_WCLK_posedge,
                            BLKEN_ipd, "BLKEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_BLKEN_WCLK_noedge_posedge,
                            tsetup_BLKEN_WCLK_noedge_posedge,
                            thold_BLKEN_WCLK_noedge_posedge,
                            thold_BLKEN_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WRAD high or low before WCLK rising
      --   Hold  WRAD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WRAD4_WCLK_posedge,
                            TmDt_WRAD4_WCLK_posedge,
                            WRAD4_ipd, "WRAD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD4_WCLK_noedge_posedge,
                            tsetup_WRAD4_WCLK_noedge_posedge,
                            thold_WRAD4_WCLK_noedge_posedge,
                            thold_WRAD4_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD3_WCLK_posedge,
                            TmDt_WRAD3_WCLK_posedge,
                            WRAD3_ipd, "WRAD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD3_WCLK_noedge_posedge,
                            tsetup_WRAD3_WCLK_noedge_posedge,
                            thold_WRAD3_WCLK_noedge_posedge,
                            thold_WRAD3_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD2_WCLK_posedge,
                            TmDt_WRAD2_WCLK_posedge,
                            WRAD2_ipd, "WRAD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD2_WCLK_noedge_posedge,
                            tsetup_WRAD2_WCLK_noedge_posedge,
                            thold_WRAD2_WCLK_noedge_posedge,
                            thold_WRAD2_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD1_WCLK_posedge,
                            TmDt_WRAD1_WCLK_posedge,
                            WRAD1_ipd, "WRAD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD1_WCLK_noedge_posedge,
                            tsetup_WRAD1_WCLK_noedge_posedge,
                            thold_WRAD1_WCLK_noedge_posedge,
                            thold_WRAD1_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      VitalSetupHoldCheck ( Tviol_WRAD0_WCLK_posedge,
                            TmDt_WRAD0_WCLK_posedge,
                            WRAD0_ipd, "WRAD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WRAD0_WCLK_noedge_posedge,
                            tsetup_WRAD0_WCLK_noedge_posedge,
                            thold_WRAD0_WCLK_noedge_posedge,
                            thold_WRAD0_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
                            
      --   Setup WD high or low before WCLK rising
      --   Hold  WD high or low before WCLK rising

      VitalSetupHoldCheck ( Tviol_WD7_WCLK_posedge,
                            TmDt_WD7_WCLK_posedge,
                            WD7_ipd, "WD7",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD7_WCLK_noedge_posedge,
                            tsetup_WD7_WCLK_noedge_posedge,
                            thold_WD7_WCLK_noedge_posedge,
                            thold_WD7_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD6_WCLK_posedge,
                            TmDt_WD6_WCLK_posedge,
                            WD6_ipd, "WD6",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD6_WCLK_noedge_posedge,
                            tsetup_WD6_WCLK_noedge_posedge,
                            thold_WD6_WCLK_noedge_posedge,
                            thold_WD6_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD5_WCLK_posedge,
                            TmDt_WD5_WCLK_posedge,
                            WD5_ipd, "WD5",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD5_WCLK_noedge_posedge,
                            tsetup_WD5_WCLK_noedge_posedge,
                            thold_WD5_WCLK_noedge_posedge,
                            thold_WD5_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD4_WCLK_posedge,
                            TmDt_WD4_WCLK_posedge,
                            WD4_ipd, "WD4",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD4_WCLK_noedge_posedge,
                            tsetup_WD4_WCLK_noedge_posedge,
                            thold_WD4_WCLK_noedge_posedge,
                            thold_WD4_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD3_WCLK_posedge,
                            TmDt_WD3_WCLK_posedge,
                            WD3_ipd, "WD3",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD3_WCLK_noedge_posedge,
                            tsetup_WD3_WCLK_noedge_posedge,
                            thold_WD3_WCLK_noedge_posedge,
                            thold_WD3_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD2_WCLK_posedge,
                            TmDt_WD2_WCLK_posedge,
                            WD2_ipd, "WD2",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD2_WCLK_noedge_posedge,
                            tsetup_WD2_WCLK_noedge_posedge,
                            thold_WD2_WCLK_noedge_posedge,
                            thold_WD2_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD1_WCLK_posedge,
                            TmDt_WD1_WCLK_posedge,
                            WD1_ipd, "WD1",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD1_WCLK_noedge_posedge,
                            tsetup_WD1_WCLK_noedge_posedge,
                            thold_WD1_WCLK_noedge_posedge,
                            thold_WD1_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      VitalSetupHoldCheck ( Tviol_WD0_WCLK_posedge,
                            TmDt_WD0_WCLK_posedge,
                            WD0_ipd, "WD0",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WD0_WCLK_noedge_posedge,
                            tsetup_WD0_WCLK_noedge_posedge,
                            thold_WD0_WCLK_noedge_posedge,
                            thold_WD0_WCLK_noedge_posedge,
                            ((To_X01(BLKEN_ipd)=BLKENS) and (To_X01(WEN_ipd)='1')),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Setup WEN high before WCLK rising
      --   Hold  WEN high after WCLK rising

      VitalSetupHoldCheck ( Tviol_WEN_WCLK_posedge,
                            TmDt_WEN_WCLK_posedge,
                            WEN_ipd, "WEN",
                            0.0 ns,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
                            tsetup_WEN_WCLK_noedge_posedge,
                            tsetup_WEN_WCLK_noedge_posedge,
                            thold_WEN_WCLK_noedge_posedge,
                            thold_WEN_WCLK_noedge_posedge,
                            (To_X01(BLKEN_ipd)=BLKENS),
                            '/',
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );

      --   Period of WCLK 

      VitalPeriodPulseCheck ( Pviol_WCLK,
                            PeriodData_WCLK,
                            WCLK_ipd, "WCLK",
                            0.0 ns,
			    tpw_WCLK_posedge + tpw_WCLK_negedge,
                            tpw_WCLK_posedge,
                            tpw_WCLK_negedge,
                            TimingCheckOn,
                            InstancePath & "/RAM8RR",
                            TRUE,
                            TRUE,
                            ERROR
                            );
    
    end if;
    
      -- #########################################################
      -- # Write Functional Section
      -- #########################################################

      -- Convert Write Address Signal to Integer
      WADDR := ((INT(WRAD4_delayed)*16)+(INT(WRAD3_delayed)*8)+(INT(WRAD2_delayed)*4)
		+(INT(WRAD1_delayed)*2)+(INT(WRAD0_delayed)));

      if (TO_X01(WCLK_ipd)='X') then
        if (TO_X01(WCLK_previous) /= 'X') then
	  assert false
	  report ": WCLK unknown"
	  severity Warning;
	end if;
      elsif (WCLK_ipd'event and (TO_X01(WCLK_ipd)='1')) then
	case TO_X01(WEN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (TO_X01(BLKEN_delayed) = 'X') then
              if (TO_X01(BLKEN_previous) /= 'X') then
	        assert false
	        report ": BLKEN unknown"
	        severity Warning;
	      end if;
	    elsif (TO_X01(BLKEN_delayed) = BLKENS) then
	      if (WADDR < 0) then
		if (TO_X01(WRAD4_delayed) = 'X') and (TO_X01(WRAD4_previous) /= 'X') then
		  assert false
		  report ": WRAD4 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD3_delayed) = 'X') and (TO_X01(WRAD3_previous) /= 'X') then
		  assert false
		  report ": WRAD3 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD2_delayed) = 'X') and (TO_X01(WRAD2_previous) /= 'X') then
		  assert false
		  report ": WRAD2 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD1_delayed) = 'X') and (TO_X01(WRAD1_previous) /= 'X') then
		  assert false
		  report ": WRAD1 unknown"
		  severity Warning;
		end if;
		if (TO_X01(WRAD0_delayed) = 'X') and (TO_X01(WRAD0_previous) /= 'X') then
		  assert false
		  report ": WRAD0 unknown"
		  severity Warning;
		end if;
	      else 
		RAM_TMP(WADDR) <= WD7_delayed & WD6_delayed & WD5_delayed & 
                                  WD4_delayed & WD3_delayed & WD2_delayed &
                                  WD1_delayed & WD0_delayed ; 
	      end if;
	    else
	      null;
	    end if;
	  when others =>
            if (TO_X01(WEN_previous) /= 'X') then
	      assert false
	      report ": WEN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;

      -- #########################################################
      -- # Read Functional Section
      -- #########################################################

      -- Convert Read Address Signal to Integer
      RADDR := ((INT(RDAD4_delayed)*16)+(INT(RDAD3_delayed)*8)+(INT(RDAD2_delayed)*4)
		+(INT(RDAD1_delayed)*2)+(INT(RDAD0_delayed)));

      if (TO_X01(RCLK_ipd) = 'X') then
	RD7_zd := 'X';
	RD6_zd := 'X';
	RD5_zd := 'X';
	RD4_zd := 'X';
	RD3_zd := 'X';
	RD2_zd := 'X';
	RD1_zd := 'X';
	RD0_zd := 'X';
	if (TO_X01(RCLK_previous) /= 'X') then
	  assert false
	  report ": RCLK unknown"
	  severity Warning;
	end if;
      elsif (RCLK_ipd'event and (TO_X01(RCLK_ipd) = '1')) then
	case TO_X01(REN_delayed) is
	  when '0' =>
	    null;
	  when '1' =>
	    if (RADDR < 0) then
	      RD7_zd := 'X';
	      RD6_zd := 'X';
	      RD5_zd := 'X';
	      RD4_zd := 'X';
	      RD3_zd := 'X';
	      RD2_zd := 'X';
	      RD1_zd := 'X';
	      RD0_zd := 'X';
	      if (TO_X01(RDAD4_delayed) = 'X') and (TO_X01(RDAD4_previous) /= 'X') then
		assert false
		report ": RDAD4 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD3_delayed) = 'X') and (TO_X01(RDAD3_previous) /= 'X') then
		assert false
		report ": RDAD3 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD2_delayed) = 'X') and (TO_X01(RDAD2_previous) /= 'X') then
		assert false
		report ": RDAD2 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD1_delayed) = 'X') and (TO_X01(RDAD1_previous) /= 'X') then
		assert false
		report ": RDAD1 unknown"
		severity Warning;
	      end if;
	      if (TO_X01(RDAD0_delayed) = 'X') and (TO_X01(RDAD0_previous) /= 'X') then
		assert false
		report ": RDAD0 unknown"
		severity Warning;
	      end if;
	    else
	      RD7_zd := RAM_TMP(RADDR)(7);
	      RD6_zd := RAM_TMP(RADDR)(6);
	      RD5_zd := RAM_TMP(RADDR)(5);
	      RD4_zd := RAM_TMP(RADDR)(4);
	      RD3_zd := RAM_TMP(RADDR)(3);
	      RD2_zd := RAM_TMP(RADDR)(2);
	      RD1_zd := RAM_TMP(RADDR)(1);
	      RD0_zd := RAM_TMP(RADDR)(0);
	    end if;
	  when others =>
	    RD7_zd := 'X';
	    RD6_zd := 'X';
	    RD5_zd := 'X';
	    RD4_zd := 'X';
	    RD3_zd := 'X';
	    RD2_zd := 'X';
	    RD1_zd := 'X';
	    RD0_zd := 'X';
            if (TO_X01(REN_previous) /= 'X') then
	      assert false
	      report ": REN unknown"
	      severity Warning;
	    end if;
	end case;
      end if;
      
      WCLK_previous := WCLK_ipd;
      RCLK_previous := RCLK_ipd;
      WEN_previous := WEN_delayed;
      REN_previous := REN_delayed;
      WEN_delayed := WEN_ipd;
      REN_delayed := REN_ipd;
      BLKEN_previous := BLKEN_delayed;
      BLKEN_delayed := BLKEN_ipd;
      WD7_delayed := WD7_ipd;
      WD6_delayed := WD6_ipd;
      WD5_delayed := WD5_ipd;
      WD4_delayed := WD4_ipd;
      WD3_delayed := WD3_ipd;
      WD2_delayed := WD2_ipd;
      WD1_delayed := WD1_ipd;
      WD0_delayed := WD0_ipd;
      WRAD4_previous := WRAD4_delayed;
      WRAD3_previous := WRAD3_delayed;
      WRAD2_previous := WRAD2_delayed;
      WRAD1_previous := WRAD1_delayed;
      WRAD0_previous := WRAD0_delayed;
      WRAD4_delayed := WRAD4_ipd;
      WRAD3_delayed := WRAD3_ipd;
      WRAD2_delayed := WRAD2_ipd;
      WRAD1_delayed := WRAD1_ipd;
      WRAD0_delayed := WRAD0_ipd;
      RDAD4_previous := RDAD4_delayed;
      RDAD3_previous := RDAD3_delayed;
      RDAD2_previous := RDAD2_delayed;
      RDAD1_previous := RDAD1_delayed;
      RDAD0_previous := RDAD0_delayed;
      RDAD4_delayed := RDAD4_ipd;
      RDAD3_delayed := RDAD3_ipd;
      RDAD2_delayed := RDAD2_ipd;
      RDAD1_delayed := RDAD1_ipd;
      RDAD0_delayed := RDAD0_ipd;

    -- #########################################################
    -- # Path Delay Section 
    -- #########################################################

    VitalPathDelay01Z (
	OutSignal => RD7,
	GlitchData => RD7_GlitchData,
	OutSignalName => "RD7",
	OutTemp => RD7_zd,
	Paths => (0 => (RCLK_ipd'last_event, 
			VitalExtendToFillDelay(tpd_RCLK_RD7), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD6,
	GlitchData => RD6_GlitchData,
	OutSignalName => "RD6",
	OutTemp => RD6_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD6), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD5,
	GlitchData => RD5_GlitchData,
	OutSignalName => "RD5",
	OutTemp => RD5_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD5), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD4,
	GlitchData => RD4_GlitchData,
	OutSignalName => "RD4",
	OutTemp => RD4_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD4), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD3,
	GlitchData => RD3_GlitchData,
	OutSignalName => "RD3",
	OutTemp => RD3_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD3), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD2,
	GlitchData => RD2_GlitchData,
	OutSignalName => "RD2",
	OutTemp => RD2_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD2), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD1,
	GlitchData => RD1_GlitchData,
	OutSignalName => "RD1",
	OutTemp => RD1_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD1), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

    VitalPathDelay01Z (
	OutSignal => RD0,
	GlitchData => RD0_GlitchData,
	OutSignalName => "RD0",
	OutTemp => RD0_zd,
	Paths => (0 => (RCLK_ipd'last_event,
			VitalExtendToFillDelay(tpd_RCLK_RD0), TRUE)
		 ),
	DefaultDelay => VitalZeroDelay01Z,
	Mode => Onevent,
	XON => TRUE,
	MsgOn => TRUE,
	MsgSeverity => WARNING
	);

  end process VITALBehavior;

end VITAL_ACT;
----- CELL TBDLHS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TBDLHS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_G_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      thold_D_G_noedge_negedge                      :	VitalDelayType := 0.000 ns;
      tsetup_D_G_noedge_negedge                     :	VitalDelayType := 0.000 ns;
      tpw_G_posedge                  :	VitalDelayType := 0.000 ns;
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_G                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      G                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TBDLHS : entity is TRUE;
end TBDLHS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of TBDLHS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';
   SIGNAL G_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   VitalWireDelay (G_ipd, G, tipd_G);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd, G_ipd)

   -- timing check results
   VARIABLE Tviol_D_G_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_D_G_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_G	: STD_ULOGIC := '0';
   VARIABLE PInfo_G	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_PAD : STD_LOGIC_VECTOR(0 to 1);
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zdi : STD_LOGIC is Results(1);
   VARIABLE PAD_zd : STD_ULOGIC := 'X';

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_D_G_negedge,
          TimingData              => Tmkr_D_G_negedge,
          TestSignal              => D_ipd,
          TestSignalName          => "D",
          TestDelay               => 0 ns,
          RefSignal               => G_ipd,
          RefSignalName          => "G",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_D_G_noedge_negedge,
          SetupLow                => tsetup_D_G_noedge_negedge,
          HoldHigh                => thold_D_G_noedge_negedge,
          HoldLow                 => thold_D_G_noedge_negedge,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/TBDLHS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_G,
          PeriodData              => PInfo_G,
          TestSignal              => G_ipd,
          TestSignalName          => "G",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => tpw_G_posedge,
          PulseWidthLow           => 0 ns,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TBDLHS",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_D_G_negedge or Pviol_G;
      VitalStateTable(
        Result => PAD_zdi,
        PreviousDataIn => PrevData_PAD,
        StateTable => DL1_Q_tab,
        DataIn => (
               D_ipd, G_ipd));
      PAD_zdi := Violation XOR PAD_zdi;
      PAD_zd := VitalBUFIF0 (data => PAD_zdi,
             enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE),
                 1 => (G_ipd'last_event, VitalExtendToFillDelay(tpd_G_PAD), TRUE),
                 2 => (E_ipd'last_event, tpd_E_PAD, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_TBDLHS_VITAL of TBDLHS is
   for VITAL_ACT
   end for;
end CFG_TBDLHS_VITAL;


----- CELL TBHS -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TBHS is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TBHS : entity is TRUE;
end TBHS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of TBHS is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_PAD, TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_TBHS_VITAL of TBHS is
   for VITAL_ACT
   end for;
end CFG_TBHS_VITAL;


----- CELL TF1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TF1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_T_CLK_noedge_posedge                    :	VitalDelayType := 0.000 ns;
      tsetup_T_CLK_noedge_posedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_posedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_posedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_posedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TF1A : entity is TRUE;
end TF1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of TF1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL T_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (T_ipd, T, tipd_T);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (T_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_T_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_posedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_posedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT TF1A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  H,  x,  H ),
    ( H,  L,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  H,  x,  L ),
    ( x,  L,  H,  H,  H,  x,  L ),
    ( U,  x,  x,  L,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_T_CLK_posedge,
          TimingData              => Tmkr_T_CLK_posedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_T_CLK_noedge_posedge,
          SetupLow                => tsetup_T_CLK_noedge_posedge,
          HoldHigh                => thold_T_CLK_noedge_posedge,
          HoldLow                 => thold_T_CLK_noedge_posedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TF1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_posedge,
          TimingData              => Tmkr_CLR_CLK_posedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_posedge,
          Removal                 => thold_CLR_CLK_noedge_posedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'R',
          HeaderMsg               => InstancePath & "/TF1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_posedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TF1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TF1A",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_T_CLK_posedge or Tviol_CLR_CLK_posedge or Pviol_CLK or Pviol_CLR;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TF1A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_delayed, T_delayed, Q_zd, CLK_ipd));
      Q_zd := Violation XOR Q_zd;
      T_delayed := T_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_TF1A_VITAL of TF1A is
   for VITAL_ACT
   end for;
end CFG_TF1A_VITAL;


----- CELL TF1B -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TF1B is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_CLR_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_CLK_Q                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      thold_T_CLK_noedge_negedge                    :	VitalDelayType := 0.000 ns;
      tsetup_T_CLK_noedge_negedge                   :	VitalDelayType := 0.000 ns;
      thold_CLR_CLK_noedge_negedge                  :	VitalDelayType := 0.000 ns;
      trecovery_CLR_CLK_posedge_negedge              :	VitalDelayType := 0.000 ns;
      tperiod_CLK_negedge            :	VitalDelayType := 0.000 ns;
      tpw_CLK_posedge                :	VitalDelayType := 0.000 ns;
      tpw_CLK_negedge                :	VitalDelayType := 0.000 ns;
      tpw_CLR_negedge                :	VitalDelayType := 0.000 ns;
      tipd_T                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLK                       :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_CLR                       :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      T                              :	in    STD_ULOGIC;
      CLK                            :	in    STD_ULOGIC;
      CLR                            :	in    STD_ULOGIC;
      Q                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TF1B : entity is TRUE;
end TF1B;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of TF1B is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL T_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLK_ipd	 : STD_ULOGIC := 'X';
   SIGNAL CLR_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (T_ipd, T, tipd_T);
   VitalWireDelay (CLK_ipd, CLK, tipd_CLK);
   VitalWireDelay (CLR_ipd, CLR, tipd_CLR);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (T_ipd, CLK_ipd, CLR_ipd)

   -- timing check results
   VARIABLE Tviol_T_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_T_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Tviol_CLR_CLK_negedge	: STD_ULOGIC := '0';
   VARIABLE Tmkr_CLR_CLK_negedge	: VitalTimingDataType := VitalTimingDataInit;
   VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
   VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
   VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

   -- functionality results
   VARIABLE Violation : STD_ULOGIC := '0';
   VARIABLE PrevData_Q : STD_LOGIC_VECTOR(0 to 4);
   VARIABLE T_delayed : STD_ULOGIC := 'X';
   VARIABLE CLK_delayed : STD_ULOGIC := 'X';
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Q_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Q_GlitchData	: VitalGlitchDataType;

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

   CONSTANT TF1A_Q_tab : VitalStateTableType := (
    ( L,  x,  x,  x,  x,  x,  L ),
    ( H,  L,  L,  H,  H,  x,  H ),
    ( H,  L,  H,  L,  H,  x,  H ),
    ( H,  H,  x,  x,  x,  x,  S ),
    ( H,  x,  x,  x,  L,  x,  S ),
    ( x,  L,  L,  L,  H,  x,  L ),
    ( x,  L,  H,  H,  H,  x,  L ),
    ( U,  x,  x,  L,  x,  x,  L ));

   begin

      ------------------------
      --  Timing Check Section
      ------------------------
      if (TimingChecksOn) then
         VitalSetupHoldCheck (
          Violation               => Tviol_T_CLK_negedge,
          TimingData              => Tmkr_T_CLK_negedge,
          TestSignal              => T_ipd,
          TestSignalName          => "T",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          SetupHigh               => tsetup_T_CLK_noedge_negedge,
          SetupLow                => tsetup_T_CLK_noedge_negedge,
          HoldHigh                => thold_T_CLK_noedge_negedge,
          HoldLow                 => thold_T_CLK_noedge_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/TF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalRecoveryRemovalCheck (
          Violation               => Tviol_CLR_CLK_negedge,
          TimingData              => Tmkr_CLR_CLK_negedge,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          RefSignal               => CLK_ipd,
          RefSignalName          => "CLK",
          RefDelay                => 0 ns,
          Recovery                => trecovery_CLR_CLK_posedge_negedge,
          Removal                 => thold_CLR_CLK_noedge_negedge,
          ActiveLow               => TRUE,
          CheckEnabled            => 
                           TRUE,
          RefTransition           => 'F',
          HeaderMsg               => InstancePath & "/TF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLK,
          PeriodData              => PInfo_CLK,
          TestSignal              => CLK_ipd,
          TestSignalName          => "CLK",
          TestDelay               => 0 ns,
          Period                  => tperiod_CLK_negedge,
          PulseWidthHigh          => tpw_CLK_posedge,
          PulseWidthLow           => tpw_CLK_negedge,
          CheckEnabled            => 
                           TO_X01((NOT CLR_ipd) ) /= '1',
          HeaderMsg               => InstancePath &"/TF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
         VitalPeriodPulseCheck (
          Violation               => Pviol_CLR,
          PeriodData              => PInfo_CLR,
          TestSignal              => CLR_ipd,
          TestSignalName          => "CLR",
          TestDelay               => 0 ns,
          Period                  => 0 ns,
          PulseWidthHigh          => 0 ns,
          PulseWidthLow           => tpw_CLR_negedge,
          CheckEnabled            => 
                           TRUE,
          HeaderMsg               => InstancePath &"/TF1B",
          Xon                     => Xon,
          MsgOn                   => MsgOn,
          MsgSeverity             => WARNING);
      end if;

      -------------------------
      --  Functionality Section
      -------------------------
      Violation := Tviol_T_CLK_negedge or Tviol_CLR_CLK_negedge or Pviol_CLR or Pviol_CLK;
      VitalStateTable(
        Result => Q_zd,
        PreviousDataIn => PrevData_Q,
        StateTable => TF1A_Q_tab,
        DataIn => (
               CLR_ipd, CLK_ipd, T_delayed, Q_zd, CLK_delayed));
      Q_zd := Violation XOR Q_zd;
      T_delayed := T_ipd;
      CLK_delayed := CLK_ipd;

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Q,
       GlitchData => Q_GlitchData,
       OutSignalName => "Q",
       OutTemp => Q_zd,
       Paths => (0 => (CLR_ipd'last_event, tpd_CLR_Q, TRUE),
                 1 => (CLK_ipd'last_event, tpd_CLK_Q, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_TF1B_VITAL of TF1B is
   for VITAL_ACT
   end for;
end CFG_TF1B_VITAL;


----- CELL TRIBUFF -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity TRIBUFF is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_E_PAD                      :	VitalDelayType01z := 
               (0.000 ns, 0.000 ns, 1.000 ns, 1.000 ns, 1.000 ns, 1.000 ns);
      tpd_D_PAD                      :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_D                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_E                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      D                              :	in    STD_ULOGIC;
      E                              :	in    STD_ULOGIC;
      PAD                            :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of TRIBUFF : entity is TRUE;
end TRIBUFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of TRIBUFF is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL D_ipd	 : STD_ULOGIC := 'X';
   SIGNAL E_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (D_ipd, D, tipd_D);
   VitalWireDelay (E_ipd, E, tipd_E);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, E_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS PAD_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE PAD_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      PAD_zd := VitalBUFIF0 (data => D_ipd,
              enable => (NOT E_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01Z (
       OutSignal => PAD,
       GlitchData => PAD_GlitchData,
       OutSignalName => "PAD",
       OutTemp => PAD_zd,
       Paths => (0 => (E_ipd'last_event, tpd_E_PAD, TRUE),
                 1 => (D_ipd'last_event, VitalExtendToFillDelay(tpd_D_PAD), TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING,
       OutputMap => "UX01ZWLH-");

end process;

end VITAL_ACT;

configuration CFG_TRIBUFF_VITAL of TRIBUFF is
   for VITAL_ACT
   end for;
end CFG_TRIBUFF_VITAL;


----- CELL VCC -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity VCC is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True);

   port(
      Y                              :	out   STD_ULOGIC := '1');
attribute VITAL_LEVEL0 of VCC : entity is TRUE;
end VCC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of VCC is
   attribute VITAL_LEVEL0 of VITAL_ACT : architecture is TRUE;


begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   --  empty
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   Y <= '1';



end VITAL_ACT;

configuration CFG_VCC_VITAL of VCC is
   for VITAL_ACT
   end for;
end CFG_VCC_VITAL;



----- CELL XA1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XA1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XA1 : entity is TRUE;
end XA1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of XA1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) AND ((B_ipd) XOR (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_XA1_VITAL of XA1 is
   for VITAL_ACT
   end for;
end CFG_XA1_VITAL;


----- CELL XA1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XA1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XA1A : entity is TRUE;
end XA1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of XA1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) AND ((NOT ((B_ipd) XOR (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_XA1A_VITAL of XA1A is
   for VITAL_ACT
   end for;
end CFG_XA1A_VITAL;


----- CELL XNOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XNOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XNOR2 : entity is TRUE;
end XNOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of XNOR2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (NOT ((B_ipd) XOR (A_ipd)));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_XNOR2_VITAL of XNOR2 is
   for VITAL_ACT
   end for;
end CFG_XNOR2_VITAL;


----- CELL XO1 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XO1 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XO1 : entity is TRUE;
end XO1;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of XO1 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR ((B_ipd) XOR (A_ipd));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_XO1_VITAL of XO1 is
   for VITAL_ACT
   end for;
end CFG_XO1_VITAL;


----- CELL XO1A -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XO1A is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_C_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_C                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      C                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XO1A : entity is TRUE;
end XO1A;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of XO1A is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';
   SIGNAL C_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   VitalWireDelay (C_ipd, C, tipd_C);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd, C_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (C_ipd) OR ((NOT ((B_ipd) XOR (A_ipd))));

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE),
                 2 => (C_ipd'last_event, tpd_C_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_XO1A_VITAL of XO1A is
   for VITAL_ACT
   end for;
end CFG_XO1A_VITAL;


----- CELL XOR2 -----
library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;


-- entity declaration --
entity XOR2 is
   generic(
      TimingChecksOn: Boolean := True;
      InstancePath: STRING := "*";
      Xon: Boolean := False;
      MsgOn: Boolean := True;
      tpd_B_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tpd_A_Y                        :	VitalDelayType01 := (1.000 ns, 1.000 ns);
      tipd_A                         :	VitalDelayType01 := (0.000 ns, 0.000 ns);
      tipd_B                         :	VitalDelayType01 := (0.000 ns, 0.000 ns));

   port(
      A                              :	in    STD_ULOGIC;
      B                              :	in    STD_ULOGIC;
      Y                              :	out   STD_ULOGIC);
attribute VITAL_LEVEL0 of XOR2 : entity is TRUE;
end XOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a42mx;
use a42mx.VTABLES.all;
architecture VITAL_ACT of XOR2 is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is TRUE;

   SIGNAL A_ipd	 : STD_ULOGIC := 'X';
   SIGNAL B_ipd	 : STD_ULOGIC := 'X';

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block
   begin
   VitalWireDelay (A_ipd, A, tipd_A);
   VitalWireDelay (B_ipd, B, tipd_B);
   end block;
   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (A_ipd, B_ipd)


   -- functionality results
   VARIABLE Results : STD_LOGIC_VECTOR(1 to 1) := (others => 'X');
   ALIAS Y_zd : STD_LOGIC is Results(1);

   -- output glitch detection variables
   VARIABLE Y_GlitchData	: VitalGlitchDataType;

   begin

      -------------------------
      --  Functionality Section
      -------------------------
      Y_zd := (B_ipd) XOR (A_ipd);

      ----------------------
      --  Path Delay Section
      ----------------------
      VitalPathDelay01 (
       OutSignal => Y,
       GlitchData => Y_GlitchData,
       OutSignalName => "Y",
       OutTemp => Y_zd,
       Paths => (0 => (B_ipd'last_event, tpd_B_Y, TRUE),
                 1 => (A_ipd'last_event, tpd_A_Y, TRUE)),
       Mode => OnDetect,
       Xon => Xon,
       MsgOn => MsgOn,
       MsgSeverity => WARNING);

end process;

end VITAL_ACT;

configuration CFG_XOR2_VITAL of XOR2 is
   for VITAL_ACT
   end for;
end CFG_XOR2_VITAL;


---- end of library ----
