*DPST Relay Subcircuit Parameters
*PULLIN     = Pull in voltage
*DROPOFF    = Drop off voltage
*CONTACT    = Contact resistance
*RESISTANCE = Coil resistance
*INDUCTANCE = Coil Inductance 
* jjt 15/6/2002: changed DPDT model to DPST.
*
*Generic DPST Relay
*Connections:     NO_A1
*                 | NO_A2
*                 | | NO_B1
*                 | | | NO_B2
*                 | | | |  T1
*                 | | | |  | T2
*                 | | | |  | |
*                 | | | |  | |
*                 | | | |  | |
*                 | | | |  | |
.SUBCKT DPSTRELAY 1 2 3 10 4 5
+ PARAMS: PULLIN=4 DROPOFF=0.1 CONTACT=1m RESISTANCE=500 INDUCTANCE=10m
L1 4 6 {(INDUCTANCE/2)}
L2 5 7 {(INDUCTANCE/2)}
R1 6 7 {RESISTANCE}
*
BNO1 8 0 V={PULLIN}-abs(v(6,7))
SW1 1 2 8 0 SWNO OFF
*
BNO2 9 0 V={PULLIN}-abs(v(6,7))
SW2 3 10 9 0 SWNO OFF
*
.MODEL SWNO SW(VT={(PULLIN*0.98)} RON={CONTACT} )
.ENDS DPSTRELAY