///////////////////////////////////////////////////////////
//  Copyright (c) 1995/2006 Xilinx Inc.
//  All Right Reserved.
///////////////////////////////////////////////////////////
//
//   ____   ___
//  /   /\/   / 
// /___/  \  /    Vendor      : Xilinx 
// \  \    \/     Version     : 8.2i 
//  \  \          Description : 
//  /  /                      
// /__/   /\      Filename    : X_PPC440.v
// \  \  /  \     Timestamp   : Fri Apr 20 13:25:10 2007

//  \__\/\__ \                    
//                                 
//  Generated by : SmartModelVerilogFileWriter (sm_verilog)
//  Revision:
///////////////////////////////////////////////////////////

`timescale 1 ps / 1 ps 

module X_PPC440 (
	APUFCMDECFPUOP,
	APUFCMDECLDSTXFERSIZE,
	APUFCMDECLOAD,
	APUFCMDECNONAUTON,
	APUFCMDECSTORE,
	APUFCMDECUDI,
	APUFCMDECUDIVALID,
	APUFCMENDIAN,
	APUFCMFLUSH,
	APUFCMINSTRUCTION,
	APUFCMINSTRVALID,
	APUFCMLOADBYTEADDR,
	APUFCMLOADDATA,
	APUFCMLOADDVALID,
	APUFCMMSRFE0,
	APUFCMMSRFE1,
	APUFCMNEXTINSTRREADY,
	APUFCMOPERANDVALID,
	APUFCMRADATA,
	APUFCMRBDATA,
	APUFCMWRITEBACKOK,
	C440CPMCORESLEEPREQ,
	C440CPMDECIRPTREQ,
	C440CPMFITIRPTREQ,
	C440CPMMSRCE,
	C440CPMMSREE,
	C440CPMTIMERRESETREQ,
	C440CPMWDIRPTREQ,
	C440DBGSYSTEMCONTROL,
	C440JTGTDO,
	C440JTGTDOEN,
	C440MACHINECHECK,
	C440RSTCHIPRESETREQ,
	C440RSTCORERESETREQ,
	C440RSTSYSTEMRESETREQ,
	C440TRCBRANCHSTATUS,
	C440TRCCYCLE,
	C440TRCEXECUTIONSTATUS,
	C440TRCTRACESTATUS,
	C440TRCTRIGGEREVENTOUT,
	C440TRCTRIGGEREVENTTYPE,
	DMA0LLRSTENGINEACK,
	DMA0LLRXDSTRDYN,
	DMA0LLTXD,
	DMA0LLTXEOFN,
	DMA0LLTXEOPN,
	DMA0LLTXREM,
	DMA0LLTXSOFN,
	DMA0LLTXSOPN,
	DMA0LLTXSRCRDYN,
	DMA0RXIRQ,
	DMA0TXIRQ,
	DMA1LLRSTENGINEACK,
	DMA1LLRXDSTRDYN,
	DMA1LLTXD,
	DMA1LLTXEOFN,
	DMA1LLTXEOPN,
	DMA1LLTXREM,
	DMA1LLTXSOFN,
	DMA1LLTXSOPN,
	DMA1LLTXSRCRDYN,
	DMA1RXIRQ,
	DMA1TXIRQ,
	DMA2LLRSTENGINEACK,
	DMA2LLRXDSTRDYN,
	DMA2LLTXD,
	DMA2LLTXEOFN,
	DMA2LLTXEOPN,
	DMA2LLTXREM,
	DMA2LLTXSOFN,
	DMA2LLTXSOPN,
	DMA2LLTXSRCRDYN,
	DMA2RXIRQ,
	DMA2TXIRQ,
	DMA3LLRSTENGINEACK,
	DMA3LLRXDSTRDYN,
	DMA3LLTXD,
	DMA3LLTXEOFN,
	DMA3LLTXEOPN,
	DMA3LLTXREM,
	DMA3LLTXSOFN,
	DMA3LLTXSOPN,
	DMA3LLTXSRCRDYN,
	DMA3RXIRQ,
	DMA3TXIRQ,
	MIMCADDRESS,
	MIMCADDRESSVALID,
	MIMCBANKCONFLICT,
	MIMCBYTEENABLE,
	MIMCREADNOTWRITE,
	MIMCROWCONFLICT,
	MIMCWRITEDATA,
	MIMCWRITEDATAVALID,
	PPCCPMINTERCONNECTBUSY,
	PPCDMDCRABUS,
	PPCDMDCRDBUSOUT,
	PPCDMDCRREAD,
	PPCDMDCRUABUS,
	PPCDMDCRWRITE,
	PPCDSDCRACK,
	PPCDSDCRDBUSIN,
	PPCDSDCRTIMEOUTWAIT,
	PPCEICINTERCONNECTIRQ,
	PPCMPLBABORT,
	PPCMPLBABUS,
	PPCMPLBBE,
	PPCMPLBBUSLOCK,
	PPCMPLBLOCKERR,
	PPCMPLBPRIORITY,
	PPCMPLBRDBURST,
	PPCMPLBREQUEST,
	PPCMPLBRNW,
	PPCMPLBSIZE,
	PPCMPLBTATTRIBUTE,
	PPCMPLBTYPE,
	PPCMPLBUABUS,
	PPCMPLBWRBURST,
	PPCMPLBWRDBUS,
	PPCS0PLBADDRACK,
	PPCS0PLBMBUSY,
	PPCS0PLBMIRQ,
	PPCS0PLBMRDERR,
	PPCS0PLBMWRERR,
	PPCS0PLBRDBTERM,
	PPCS0PLBRDCOMP,
	PPCS0PLBRDDACK,
	PPCS0PLBRDDBUS,
	PPCS0PLBRDWDADDR,
	PPCS0PLBREARBITRATE,
	PPCS0PLBSSIZE,
	PPCS0PLBWAIT,
	PPCS0PLBWRBTERM,
	PPCS0PLBWRCOMP,
	PPCS0PLBWRDACK,
	PPCS1PLBADDRACK,
	PPCS1PLBMBUSY,
	PPCS1PLBMIRQ,
	PPCS1PLBMRDERR,
	PPCS1PLBMWRERR,
	PPCS1PLBRDBTERM,
	PPCS1PLBRDCOMP,
	PPCS1PLBRDDACK,
	PPCS1PLBRDDBUS,
	PPCS1PLBRDWDADDR,
	PPCS1PLBREARBITRATE,
	PPCS1PLBSSIZE,
	PPCS1PLBWAIT,
	PPCS1PLBWRBTERM,
	PPCS1PLBWRCOMP,
	PPCS1PLBWRDACK,

	CPMC440CLK,
	CPMC440CLKEN,
	CPMC440CORECLOCKINACTIVE,
	CPMC440TIMERCLOCK,
	CPMDCRCLK,
	CPMDMA0LLCLK,
	CPMDMA1LLCLK,
	CPMDMA2LLCLK,
	CPMDMA3LLCLK,
	CPMFCMCLK,
	CPMINTERCONNECTCLK,
	CPMINTERCONNECTCLKEN,
	CPMINTERCONNECTCLKNTO1,
	CPMMCCLK,
	CPMPPCMPLBCLK,
	CPMPPCS0PLBCLK,
	CPMPPCS1PLBCLK,
	DBGC440DEBUGHALT,
	DBGC440SYSTEMSTATUS,
	DBGC440UNCONDDEBUGEVENT,
	DCRPPCDMACK,
	DCRPPCDMDBUSIN,
	DCRPPCDMTIMEOUTWAIT,
	DCRPPCDSABUS,
	DCRPPCDSDBUSOUT,
	DCRPPCDSREAD,
	DCRPPCDSWRITE,
	EICC440CRITIRQ,
	EICC440EXTIRQ,
	FCMAPUCONFIRMINSTR,
	FCMAPUCR,
	FCMAPUDONE,
	FCMAPUEXCEPTION,
	FCMAPUFPSCRFEX,
	FCMAPURESULT,
	FCMAPURESULTVALID,
	FCMAPUSLEEPNOTREADY,
	FCMAPUSTOREDATA,
	JTGC440TCK,
	JTGC440TDI,
	JTGC440TMS,
	JTGC440TRSTNEG,
	LLDMA0RSTENGINEREQ,
	LLDMA0RXD,
	LLDMA0RXEOFN,
	LLDMA0RXEOPN,
	LLDMA0RXREM,
	LLDMA0RXSOFN,
	LLDMA0RXSOPN,
	LLDMA0RXSRCRDYN,
	LLDMA0TXDSTRDYN,
	LLDMA1RSTENGINEREQ,
	LLDMA1RXD,
	LLDMA1RXEOFN,
	LLDMA1RXEOPN,
	LLDMA1RXREM,
	LLDMA1RXSOFN,
	LLDMA1RXSOPN,
	LLDMA1RXSRCRDYN,
	LLDMA1TXDSTRDYN,
	LLDMA2RSTENGINEREQ,
	LLDMA2RXD,
	LLDMA2RXEOFN,
	LLDMA2RXEOPN,
	LLDMA2RXREM,
	LLDMA2RXSOFN,
	LLDMA2RXSOPN,
	LLDMA2RXSRCRDYN,
	LLDMA2TXDSTRDYN,
	LLDMA3RSTENGINEREQ,
	LLDMA3RXD,
	LLDMA3RXEOFN,
	LLDMA3RXEOPN,
	LLDMA3RXREM,
	LLDMA3RXSOFN,
	LLDMA3RXSOPN,
	LLDMA3RXSRCRDYN,
	LLDMA3TXDSTRDYN,
	MCMIADDRREADYTOACCEPT,
	MCMIREADDATA,
	MCMIREADDATAERR,
	MCMIREADDATAVALID,
	PLBPPCMADDRACK,
	PLBPPCMMBUSY,
	PLBPPCMMIRQ,
	PLBPPCMMRDERR,
	PLBPPCMMWRERR,
	PLBPPCMRDBTERM,
	PLBPPCMRDDACK,
	PLBPPCMRDDBUS,
	PLBPPCMRDPENDPRI,
	PLBPPCMRDPENDREQ,
	PLBPPCMRDWDADDR,
	PLBPPCMREARBITRATE,
	PLBPPCMREQPRI,
	PLBPPCMSSIZE,
	PLBPPCMTIMEOUT,
	PLBPPCMWRBTERM,
	PLBPPCMWRDACK,
	PLBPPCMWRPENDPRI,
	PLBPPCMWRPENDREQ,
	PLBPPCS0ABORT,
	PLBPPCS0ABUS,
	PLBPPCS0BE,
	PLBPPCS0BUSLOCK,
	PLBPPCS0LOCKERR,
	PLBPPCS0MASTERID,
	PLBPPCS0MSIZE,
	PLBPPCS0PAVALID,
	PLBPPCS0RDBURST,
	PLBPPCS0RDPENDPRI,
	PLBPPCS0RDPENDREQ,
	PLBPPCS0RDPRIM,
	PLBPPCS0REQPRI,
	PLBPPCS0RNW,
	PLBPPCS0SAVALID,
	PLBPPCS0SIZE,
	PLBPPCS0TATTRIBUTE,
	PLBPPCS0TYPE,
	PLBPPCS0UABUS,
	PLBPPCS0WRBURST,
	PLBPPCS0WRDBUS,
	PLBPPCS0WRPENDPRI,
	PLBPPCS0WRPENDREQ,
	PLBPPCS0WRPRIM,
	PLBPPCS1ABORT,
	PLBPPCS1ABUS,
	PLBPPCS1BE,
	PLBPPCS1BUSLOCK,
	PLBPPCS1LOCKERR,
	PLBPPCS1MASTERID,
	PLBPPCS1MSIZE,
	PLBPPCS1PAVALID,
	PLBPPCS1RDBURST,
	PLBPPCS1RDPENDPRI,
	PLBPPCS1RDPENDREQ,
	PLBPPCS1RDPRIM,
	PLBPPCS1REQPRI,
	PLBPPCS1RNW,
	PLBPPCS1SAVALID,
	PLBPPCS1SIZE,
	PLBPPCS1TATTRIBUTE,
	PLBPPCS1TYPE,
	PLBPPCS1UABUS,
	PLBPPCS1WRBURST,
	PLBPPCS1WRDBUS,
	PLBPPCS1WRPENDPRI,
	PLBPPCS1WRPENDREQ,
	PLBPPCS1WRPRIM,
	RSTC440RESETCHIP,
	RSTC440RESETCORE,
	RSTC440RESETSYSTEM,
	TIEC440DCURDLDCACHEPLBPRIO,
	TIEC440DCURDNONCACHEPLBPRIO,
	TIEC440DCURDTOUCHPLBPRIO,
	TIEC440DCURDURGENTPLBPRIO,
	TIEC440DCUWRFLUSHPLBPRIO,
	TIEC440DCUWRSTOREPLBPRIO,
	TIEC440DCUWRURGENTPLBPRIO,
	TIEC440ENDIANRESET,
	TIEC440ERPNRESET,
	TIEC440ICURDFETCHPLBPRIO,
	TIEC440ICURDSPECPLBPRIO,
	TIEC440ICURDTOUCHPLBPRIO,
	TIEC440PIR,
	TIEC440PVR,
	TIEC440USERRESET,
	TIEDCRBASEADDR,
	TRCC440TRACEDISABLE,
	TRCC440TRIGGEREVENTIN

);

parameter LOC = "UNPLACED";

parameter CLOCK_DELAY = "FALSE";
parameter DCR_AUTOLOCK_ENABLE = "TRUE";
parameter PPCDM_ASYNCMODE = "FALSE";
parameter PPCDS_ASYNCMODE = "FALSE";
parameter PPCS0_WIDTH_128N64 = "TRUE";
parameter PPCS1_WIDTH_128N64 = "TRUE";
parameter [0:16] APU_CONTROL = 17'h02000;
parameter [0:23] APU_UDI0 = 24'h000000;
parameter [0:23] APU_UDI1 = 24'h000000;
parameter [0:23] APU_UDI10 = 24'h000000;
parameter [0:23] APU_UDI11 = 24'h000000;
parameter [0:23] APU_UDI12 = 24'h000000;
parameter [0:23] APU_UDI13 = 24'h000000;
parameter [0:23] APU_UDI14 = 24'h000000;
parameter [0:23] APU_UDI15 = 24'h000000;
parameter [0:23] APU_UDI2 = 24'h000000;
parameter [0:23] APU_UDI3 = 24'h000000;
parameter [0:23] APU_UDI4 = 24'h000000;
parameter [0:23] APU_UDI5 = 24'h000000;
parameter [0:23] APU_UDI6 = 24'h000000;
parameter [0:23] APU_UDI7 = 24'h000000;
parameter [0:23] APU_UDI8 = 24'h000000;
parameter [0:23] APU_UDI9 = 24'h000000;
parameter [0:31] DMA0_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA0_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA1_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA1_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA2_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA2_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA3_RXCHANNELCTRL = 32'h01010000;
parameter [0:31] DMA3_TXCHANNELCTRL = 32'h01010000;
parameter [0:31] INTERCONNECT_IMASK = 32'hFFFFFFFF;
parameter [0:31] INTERCONNECT_TMPL_SEL = 32'h3FFFFFFF;
parameter [0:31] MI_ARBCONFIG = 32'h00432010;
parameter [0:31] MI_BANKCONFLICT_MASK = 32'h00000000;
parameter [0:31] MI_CONTROL = 32'h0000008F;
parameter [0:31] MI_ROWCONFLICT_MASK = 32'h00000000;
parameter [0:31] PPCM_ARBCONFIG = 32'h00432010;
parameter [0:31] PPCM_CONTROL = 32'h8000009F;
parameter [0:31] PPCM_COUNTER = 32'h00000500;
parameter [0:31] PPCS0_ADDRMAP_TMPL0 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_ADDRMAP_TMPL1 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_ADDRMAP_TMPL2 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_ADDRMAP_TMPL3 = 32'hFFFFFFFF;
parameter [0:31] PPCS0_CONTROL = 32'h8033336C;
parameter [0:31] PPCS1_ADDRMAP_TMPL0 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_ADDRMAP_TMPL1 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_ADDRMAP_TMPL2 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_ADDRMAP_TMPL3 = 32'hFFFFFFFF;
parameter [0:31] PPCS1_CONTROL = 32'h8033336C;
parameter [0:31] XBAR_ADDRMAP_TMPL0 = 32'hFFFF0000;
parameter [0:31] XBAR_ADDRMAP_TMPL1 = 32'h00000000;
parameter [0:31] XBAR_ADDRMAP_TMPL2 = 32'h00000000;
parameter [0:31] XBAR_ADDRMAP_TMPL3 = 32'h00000000;
parameter [0:7] DMA0_CONTROL = 8'h00;
parameter [0:7] DMA1_CONTROL = 8'h00;
parameter [0:7] DMA2_CONTROL = 8'h00;
parameter [0:7] DMA3_CONTROL = 8'h00;
parameter [0:9] DMA0_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA0_TXIRQTIMER = 10'h3FF;
parameter [0:9] DMA1_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA1_TXIRQTIMER = 10'h3FF;
parameter [0:9] DMA2_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA2_TXIRQTIMER = 10'h3FF;
parameter [0:9] DMA3_RXIRQTIMER = 10'h3FF;
parameter [0:9] DMA3_TXIRQTIMER = 10'h3FF;

localparam in_delay = 1;
localparam out_delay = 0;
localparam CLK_DELAY = 0;

output APUFCMDECFPUOP;
output APUFCMDECLOAD;
output APUFCMDECNONAUTON;
output APUFCMDECSTORE;
output APUFCMDECUDIVALID;
output APUFCMENDIAN;
output APUFCMFLUSH;
output APUFCMINSTRVALID;
output APUFCMLOADDVALID;
output APUFCMMSRFE0;
output APUFCMMSRFE1;
output APUFCMNEXTINSTRREADY;
output APUFCMOPERANDVALID;
output APUFCMWRITEBACKOK;
output C440CPMCORESLEEPREQ;
output C440CPMDECIRPTREQ;
output C440CPMFITIRPTREQ;
output C440CPMMSRCE;
output C440CPMMSREE;
output C440CPMTIMERRESETREQ;
output C440CPMWDIRPTREQ;
output C440JTGTDO;
output C440JTGTDOEN;
output C440MACHINECHECK;
output C440RSTCHIPRESETREQ;
output C440RSTCORERESETREQ;
output C440RSTSYSTEMRESETREQ;
output C440TRCCYCLE;
output C440TRCTRIGGEREVENTOUT;
output DMA0LLRSTENGINEACK;
output DMA0LLRXDSTRDYN;
output DMA0LLTXEOFN;
output DMA0LLTXEOPN;
output DMA0LLTXSOFN;
output DMA0LLTXSOPN;
output DMA0LLTXSRCRDYN;
output DMA0RXIRQ;
output DMA0TXIRQ;
output DMA1LLRSTENGINEACK;
output DMA1LLRXDSTRDYN;
output DMA1LLTXEOFN;
output DMA1LLTXEOPN;
output DMA1LLTXSOFN;
output DMA1LLTXSOPN;
output DMA1LLTXSRCRDYN;
output DMA1RXIRQ;
output DMA1TXIRQ;
output DMA2LLRSTENGINEACK;
output DMA2LLRXDSTRDYN;
output DMA2LLTXEOFN;
output DMA2LLTXEOPN;
output DMA2LLTXSOFN;
output DMA2LLTXSOPN;
output DMA2LLTXSRCRDYN;
output DMA2RXIRQ;
output DMA2TXIRQ;
output DMA3LLRSTENGINEACK;
output DMA3LLRXDSTRDYN;
output DMA3LLTXEOFN;
output DMA3LLTXEOPN;
output DMA3LLTXSOFN;
output DMA3LLTXSOPN;
output DMA3LLTXSRCRDYN;
output DMA3RXIRQ;
output DMA3TXIRQ;
output MIMCADDRESSVALID;
output MIMCBANKCONFLICT;
output MIMCREADNOTWRITE;
output MIMCROWCONFLICT;
output MIMCWRITEDATAVALID;
output PPCCPMINTERCONNECTBUSY;
output PPCDMDCRREAD;
output PPCDMDCRWRITE;
output PPCDSDCRACK;
output PPCDSDCRTIMEOUTWAIT;
output PPCEICINTERCONNECTIRQ;
output PPCMPLBABORT;
output PPCMPLBBUSLOCK;
output PPCMPLBLOCKERR;
output PPCMPLBRDBURST;
output PPCMPLBREQUEST;
output PPCMPLBRNW;
output PPCMPLBWRBURST;
output PPCS0PLBADDRACK;
output PPCS0PLBRDBTERM;
output PPCS0PLBRDCOMP;
output PPCS0PLBRDDACK;
output PPCS0PLBREARBITRATE;
output PPCS0PLBWAIT;
output PPCS0PLBWRBTERM;
output PPCS0PLBWRCOMP;
output PPCS0PLBWRDACK;
output PPCS1PLBADDRACK;
output PPCS1PLBRDBTERM;
output PPCS1PLBRDCOMP;
output PPCS1PLBRDDACK;
output PPCS1PLBREARBITRATE;
output PPCS1PLBWAIT;
output PPCS1PLBWRBTERM;
output PPCS1PLBWRCOMP;
output PPCS1PLBWRDACK;
output [0:127] APUFCMLOADDATA;
output [0:127] MIMCWRITEDATA;
output [0:127] PPCMPLBWRDBUS;
output [0:127] PPCS0PLBRDDBUS;
output [0:127] PPCS1PLBRDDBUS;
output [0:13] C440TRCTRIGGEREVENTTYPE;
output [0:15] MIMCBYTEENABLE;
output [0:15] PPCMPLBBE;
output [0:15] PPCMPLBTATTRIBUTE;
output [0:1] PPCMPLBPRIORITY;
output [0:1] PPCS0PLBSSIZE;
output [0:1] PPCS1PLBSSIZE;
output [0:2] APUFCMDECLDSTXFERSIZE;
output [0:2] C440TRCBRANCHSTATUS;
output [0:2] PPCMPLBTYPE;
output [0:31] APUFCMINSTRUCTION;
output [0:31] APUFCMRADATA;
output [0:31] APUFCMRBDATA;
output [0:31] DMA0LLTXD;
output [0:31] DMA1LLTXD;
output [0:31] DMA2LLTXD;
output [0:31] DMA3LLTXD;
output [0:31] PPCDMDCRDBUSOUT;
output [0:31] PPCDSDCRDBUSIN;
output [0:31] PPCMPLBABUS;
output [0:35] MIMCADDRESS;
output [0:3] APUFCMDECUDI;
output [0:3] APUFCMLOADBYTEADDR;
output [0:3] DMA0LLTXREM;
output [0:3] DMA1LLTXREM;
output [0:3] DMA2LLTXREM;
output [0:3] DMA3LLTXREM;
output [0:3] PPCMPLBSIZE;
output [0:3] PPCS0PLBMBUSY;
output [0:3] PPCS0PLBMIRQ;
output [0:3] PPCS0PLBMRDERR;
output [0:3] PPCS0PLBMWRERR;
output [0:3] PPCS0PLBRDWDADDR;
output [0:3] PPCS1PLBMBUSY;
output [0:3] PPCS1PLBMIRQ;
output [0:3] PPCS1PLBMRDERR;
output [0:3] PPCS1PLBMWRERR;
output [0:3] PPCS1PLBRDWDADDR;
output [0:4] C440TRCEXECUTIONSTATUS;
output [0:6] C440TRCTRACESTATUS;
output [0:7] C440DBGSYSTEMCONTROL;
output [0:9] PPCDMDCRABUS;
output [20:21] PPCDMDCRUABUS;
output [28:31] PPCMPLBUABUS;

input CPMC440CLK;
input CPMC440CLKEN;
input CPMC440CORECLOCKINACTIVE;
input CPMC440TIMERCLOCK;
input CPMDCRCLK;
input CPMDMA0LLCLK;
input CPMDMA1LLCLK;
input CPMDMA2LLCLK;
input CPMDMA3LLCLK;
input CPMFCMCLK;
input CPMINTERCONNECTCLK;
input CPMINTERCONNECTCLKEN;
input CPMINTERCONNECTCLKNTO1;
input CPMMCCLK;
input CPMPPCMPLBCLK;
input CPMPPCS0PLBCLK;
input CPMPPCS1PLBCLK;
input DBGC440DEBUGHALT;
input DBGC440UNCONDDEBUGEVENT;
input DCRPPCDMACK;
input DCRPPCDMTIMEOUTWAIT;
input DCRPPCDSREAD;
input DCRPPCDSWRITE;
input EICC440CRITIRQ;
input EICC440EXTIRQ;
input FCMAPUCONFIRMINSTR;
input FCMAPUDONE;
input FCMAPUEXCEPTION;
input FCMAPUFPSCRFEX;
input FCMAPURESULTVALID;
input FCMAPUSLEEPNOTREADY;
input JTGC440TCK;
input JTGC440TDI;
input JTGC440TMS;
input JTGC440TRSTNEG;
input LLDMA0RSTENGINEREQ;
input LLDMA0RXEOFN;
input LLDMA0RXEOPN;
input LLDMA0RXSOFN;
input LLDMA0RXSOPN;
input LLDMA0RXSRCRDYN;
input LLDMA0TXDSTRDYN;
input LLDMA1RSTENGINEREQ;
input LLDMA1RXEOFN;
input LLDMA1RXEOPN;
input LLDMA1RXSOFN;
input LLDMA1RXSOPN;
input LLDMA1RXSRCRDYN;
input LLDMA1TXDSTRDYN;
input LLDMA2RSTENGINEREQ;
input LLDMA2RXEOFN;
input LLDMA2RXEOPN;
input LLDMA2RXSOFN;
input LLDMA2RXSOPN;
input LLDMA2RXSRCRDYN;
input LLDMA2TXDSTRDYN;
input LLDMA3RSTENGINEREQ;
input LLDMA3RXEOFN;
input LLDMA3RXEOPN;
input LLDMA3RXSOFN;
input LLDMA3RXSOPN;
input LLDMA3RXSRCRDYN;
input LLDMA3TXDSTRDYN;
input MCMIADDRREADYTOACCEPT;
input MCMIREADDATAERR;
input MCMIREADDATAVALID;
input PLBPPCMADDRACK;
input PLBPPCMMBUSY;
input PLBPPCMMIRQ;
input PLBPPCMMRDERR;
input PLBPPCMMWRERR;
input PLBPPCMRDBTERM;
input PLBPPCMRDDACK;
input PLBPPCMRDPENDREQ;
input PLBPPCMREARBITRATE;
input PLBPPCMTIMEOUT;
input PLBPPCMWRBTERM;
input PLBPPCMWRDACK;
input PLBPPCMWRPENDREQ;
input PLBPPCS0ABORT;
input PLBPPCS0BUSLOCK;
input PLBPPCS0LOCKERR;
input PLBPPCS0PAVALID;
input PLBPPCS0RDBURST;
input PLBPPCS0RDPENDREQ;
input PLBPPCS0RDPRIM;
input PLBPPCS0RNW;
input PLBPPCS0SAVALID;
input PLBPPCS0WRBURST;
input PLBPPCS0WRPENDREQ;
input PLBPPCS0WRPRIM;
input PLBPPCS1ABORT;
input PLBPPCS1BUSLOCK;
input PLBPPCS1LOCKERR;
input PLBPPCS1PAVALID;
input PLBPPCS1RDBURST;
input PLBPPCS1RDPENDREQ;
input PLBPPCS1RDPRIM;
input PLBPPCS1RNW;
input PLBPPCS1SAVALID;
input PLBPPCS1WRBURST;
input PLBPPCS1WRPENDREQ;
input PLBPPCS1WRPRIM;
input RSTC440RESETCHIP;
input RSTC440RESETCORE;
input RSTC440RESETSYSTEM;
input TIEC440ENDIANRESET;
input TRCC440TRACEDISABLE;
input TRCC440TRIGGEREVENTIN;
input [0:127] FCMAPUSTOREDATA;
input [0:127] MCMIREADDATA;
input [0:127] PLBPPCMRDDBUS;
input [0:127] PLBPPCS0WRDBUS;
input [0:127] PLBPPCS1WRDBUS;
input [0:15] PLBPPCS0BE;
input [0:15] PLBPPCS0TATTRIBUTE;
input [0:15] PLBPPCS1BE;
input [0:15] PLBPPCS1TATTRIBUTE;
input [0:1] PLBPPCMRDPENDPRI;
input [0:1] PLBPPCMREQPRI;
input [0:1] PLBPPCMSSIZE;
input [0:1] PLBPPCMWRPENDPRI;
input [0:1] PLBPPCS0MASTERID;
input [0:1] PLBPPCS0MSIZE;
input [0:1] PLBPPCS0RDPENDPRI;
input [0:1] PLBPPCS0REQPRI;
input [0:1] PLBPPCS0WRPENDPRI;
input [0:1] PLBPPCS1MASTERID;
input [0:1] PLBPPCS1MSIZE;
input [0:1] PLBPPCS1RDPENDPRI;
input [0:1] PLBPPCS1REQPRI;
input [0:1] PLBPPCS1WRPENDPRI;
input [0:1] TIEC440DCURDLDCACHEPLBPRIO;
input [0:1] TIEC440DCURDNONCACHEPLBPRIO;
input [0:1] TIEC440DCURDTOUCHPLBPRIO;
input [0:1] TIEC440DCURDURGENTPLBPRIO;
input [0:1] TIEC440DCUWRFLUSHPLBPRIO;
input [0:1] TIEC440DCUWRSTOREPLBPRIO;
input [0:1] TIEC440DCUWRURGENTPLBPRIO;
input [0:1] TIEC440ICURDFETCHPLBPRIO;
input [0:1] TIEC440ICURDSPECPLBPRIO;
input [0:1] TIEC440ICURDTOUCHPLBPRIO;
input [0:1] TIEDCRBASEADDR;
input [0:2] PLBPPCS0TYPE;
input [0:2] PLBPPCS1TYPE;
input [0:31] DCRPPCDMDBUSIN;
input [0:31] DCRPPCDSDBUSOUT;
input [0:31] FCMAPURESULT;
input [0:31] LLDMA0RXD;
input [0:31] LLDMA1RXD;
input [0:31] LLDMA2RXD;
input [0:31] LLDMA3RXD;
input [0:31] PLBPPCS0ABUS;
input [0:31] PLBPPCS1ABUS;
input [0:3] FCMAPUCR;
input [0:3] LLDMA0RXREM;
input [0:3] LLDMA1RXREM;
input [0:3] LLDMA2RXREM;
input [0:3] LLDMA3RXREM;
input [0:3] PLBPPCMRDWDADDR;
input [0:3] PLBPPCS0SIZE;
input [0:3] PLBPPCS1SIZE;
input [0:3] TIEC440ERPNRESET;
input [0:3] TIEC440USERRESET;
input [0:4] DBGC440SYSTEMSTATUS;
input [0:9] DCRPPCDSABUS;
input [28:31] PLBPPCS0UABUS;
input [28:31] PLBPPCS1UABUS;
input [28:31] TIEC440PIR;
input [28:31] TIEC440PVR;

reg [0:4] CLOCK_DELAY_BINARY;
reg DCR_AUTOLOCK_ENABLE_BINARY;
reg PPCDM_ASYNCMODE_BINARY;
reg PPCDS_ASYNCMODE_BINARY;
reg PPCS0_WIDTH_128N64_BINARY;
reg PPCS1_WIDTH_128N64_BINARY;

tri0 GSR = glbl.GSR;
reg notifier;

wire APUFCMDECFPUOP_OUT;
wire APUFCMDECLOAD_OUT;
wire APUFCMDECNONAUTON_OUT;
wire APUFCMDECSTORE_OUT;
wire APUFCMDECUDIVALID_OUT;
wire APUFCMENDIAN_OUT;
wire APUFCMFLUSH_OUT;
wire APUFCMINSTRVALID_OUT;
wire APUFCMLOADDVALID_OUT;
wire APUFCMMSRFE0_OUT;
wire APUFCMMSRFE1_OUT;
wire APUFCMNEXTINSTRREADY_OUT;
wire APUFCMOPERANDVALID_OUT;
wire APUFCMWRITEBACKOK_OUT;
wire C440CPMCORESLEEPREQ_OUT;
wire C440CPMDECIRPTREQ_OUT;
wire C440CPMFITIRPTREQ_OUT;
wire C440CPMMSRCE_OUT;
wire C440CPMMSREE_OUT;
wire C440CPMTIMERRESETREQ_OUT;
wire C440CPMWDIRPTREQ_OUT;
wire C440JTGTDOEN_OUT;
wire C440JTGTDO_OUT;
wire C440MACHINECHECK_OUT;
wire C440RSTCHIPRESETREQ_OUT;
wire C440RSTCORERESETREQ_OUT;
wire C440RSTSYSTEMRESETREQ_OUT;
wire C440TRCCYCLE_OUT;
wire C440TRCTRIGGEREVENTOUT_OUT;
wire DMA0LLRSTENGINEACK_OUT;
wire DMA0LLRXDSTRDYN_OUT;
wire DMA0LLTXEOFN_OUT;
wire DMA0LLTXEOPN_OUT;
wire DMA0LLTXSOFN_OUT;
wire DMA0LLTXSOPN_OUT;
wire DMA0LLTXSRCRDYN_OUT;
wire DMA0RXIRQ_OUT;
wire DMA0TXIRQ_OUT;
wire DMA1LLRSTENGINEACK_OUT;
wire DMA1LLRXDSTRDYN_OUT;
wire DMA1LLTXEOFN_OUT;
wire DMA1LLTXEOPN_OUT;
wire DMA1LLTXSOFN_OUT;
wire DMA1LLTXSOPN_OUT;
wire DMA1LLTXSRCRDYN_OUT;
wire DMA1RXIRQ_OUT;
wire DMA1TXIRQ_OUT;
wire DMA2LLRSTENGINEACK_OUT;
wire DMA2LLRXDSTRDYN_OUT;
wire DMA2LLTXEOFN_OUT;
wire DMA2LLTXEOPN_OUT;
wire DMA2LLTXSOFN_OUT;
wire DMA2LLTXSOPN_OUT;
wire DMA2LLTXSRCRDYN_OUT;
wire DMA2RXIRQ_OUT;
wire DMA2TXIRQ_OUT;
wire DMA3LLRSTENGINEACK_OUT;
wire DMA3LLRXDSTRDYN_OUT;
wire DMA3LLTXEOFN_OUT;
wire DMA3LLTXEOPN_OUT;
wire DMA3LLTXSOFN_OUT;
wire DMA3LLTXSOPN_OUT;
wire DMA3LLTXSRCRDYN_OUT;
wire DMA3RXIRQ_OUT;
wire DMA3TXIRQ_OUT;
wire MIMCADDRESSVALID_OUT;
wire MIMCBANKCONFLICT_OUT;
wire MIMCREADNOTWRITE_OUT;
wire MIMCROWCONFLICT_OUT;
wire MIMCWRITEDATAVALID_OUT;
wire PPCCPMINTERCONNECTBUSY_OUT;
wire PPCDMDCRREAD_OUT;
wire PPCDMDCRWRITE_OUT;
wire PPCDSDCRACK_OUT;
wire PPCDSDCRTIMEOUTWAIT_OUT;
wire PPCEICINTERCONNECTIRQ_OUT;
wire PPCMPLBABORT_OUT;
wire PPCMPLBBUSLOCK_OUT;
wire PPCMPLBLOCKERR_OUT;
wire PPCMPLBRDBURST_OUT;
wire PPCMPLBREQUEST_OUT;
wire PPCMPLBRNW_OUT;
wire PPCMPLBWRBURST_OUT;
wire PPCS0PLBADDRACK_OUT;
wire PPCS0PLBRDBTERM_OUT;
wire PPCS0PLBRDCOMP_OUT;
wire PPCS0PLBRDDACK_OUT;
wire PPCS0PLBREARBITRATE_OUT;
wire PPCS0PLBWAIT_OUT;
wire PPCS0PLBWRBTERM_OUT;
wire PPCS0PLBWRCOMP_OUT;
wire PPCS0PLBWRDACK_OUT;
wire PPCS1PLBADDRACK_OUT;
wire PPCS1PLBRDBTERM_OUT;
wire PPCS1PLBRDCOMP_OUT;
wire PPCS1PLBRDDACK_OUT;
wire PPCS1PLBREARBITRATE_OUT;
wire PPCS1PLBWAIT_OUT;
wire PPCS1PLBWRBTERM_OUT;
wire PPCS1PLBWRCOMP_OUT;
wire PPCS1PLBWRDACK_OUT;
wire [0:127] APUFCMLOADDATA_OUT;
wire [0:127] MIMCWRITEDATA_OUT;
wire [0:127] PPCMPLBWRDBUS_OUT;
wire [0:127] PPCS0PLBRDDBUS_OUT;
wire [0:127] PPCS1PLBRDDBUS_OUT;
wire [0:13] C440TRCTRIGGEREVENTTYPE_OUT;
wire [0:15] MIMCBYTEENABLE_OUT;
wire [0:15] PPCMPLBBE_OUT;
wire [0:15] PPCMPLBTATTRIBUTE_OUT;
wire [0:1] PPCMPLBPRIORITY_OUT;
wire [0:1] PPCS0PLBSSIZE_OUT;
wire [0:1] PPCS1PLBSSIZE_OUT;
wire [0:2] APUFCMDECLDSTXFERSIZE_OUT;
wire [0:2] C440TRCBRANCHSTATUS_OUT;
wire [0:2] PPCMPLBTYPE_OUT;
wire [0:31] APUFCMINSTRUCTION_OUT;
wire [0:31] APUFCMRADATA_OUT;
wire [0:31] APUFCMRBDATA_OUT;
wire [0:31] DMA0LLTXD_OUT;
wire [0:31] DMA1LLTXD_OUT;
wire [0:31] DMA2LLTXD_OUT;
wire [0:31] DMA3LLTXD_OUT;
wire [0:31] PPCDMDCRDBUSOUT_OUT;
wire [0:31] PPCDSDCRDBUSIN_OUT;
wire [0:31] PPCMPLBABUS_OUT;
wire [0:35] MIMCADDRESS_OUT;
wire [0:3] APUFCMDECUDI_OUT;
wire [0:3] APUFCMLOADBYTEADDR_OUT;
wire [0:3] DMA0LLTXREM_OUT;
wire [0:3] DMA1LLTXREM_OUT;
wire [0:3] DMA2LLTXREM_OUT;
wire [0:3] DMA3LLTXREM_OUT;
wire [0:3] PPCMPLBSIZE_OUT;
wire [0:3] PPCS0PLBMBUSY_OUT;
wire [0:3] PPCS0PLBMIRQ_OUT;
wire [0:3] PPCS0PLBMRDERR_OUT;
wire [0:3] PPCS0PLBMWRERR_OUT;
wire [0:3] PPCS0PLBRDWDADDR_OUT;
wire [0:3] PPCS1PLBMBUSY_OUT;
wire [0:3] PPCS1PLBMIRQ_OUT;
wire [0:3] PPCS1PLBMRDERR_OUT;
wire [0:3] PPCS1PLBMWRERR_OUT;
wire [0:3] PPCS1PLBRDWDADDR_OUT;
wire [0:4] C440TRCEXECUTIONSTATUS_OUT;
wire [0:6] C440TRCTRACESTATUS_OUT;
wire [0:7] C440DBGSYSTEMCONTROL_OUT;
wire [0:9] PPCDMDCRABUS_OUT;
wire [20:21] PPCDMDCRUABUS_OUT;
wire [28:31] PPCMPLBUABUS_OUT;

wire CPMC440CLKEN_IN;
wire CPMC440CLK_IN;
wire CPMC440CORECLOCKINACTIVE_IN;
wire CPMC440TIMERCLOCK_IN;
wire CPMDCRCLK_IN;
wire CPMDMA0LLCLK_IN;
wire CPMDMA1LLCLK_IN;
wire CPMDMA2LLCLK_IN;
wire CPMDMA3LLCLK_IN;
wire CPMFCMCLK_IN;
wire CPMINTERCONNECTCLKEN_IN;
wire CPMINTERCONNECTCLKNTO1_IN;
wire CPMINTERCONNECTCLK_IN;
wire CPMMCCLK_IN;
wire CPMPPCMPLBCLK_IN;
wire CPMPPCS0PLBCLK_IN;
wire CPMPPCS1PLBCLK_IN;
wire DBGC440DEBUGHALT_IN;
wire DBGC440UNCONDDEBUGEVENT_IN;
wire DCRPPCDMACK_IN;
wire DCRPPCDMTIMEOUTWAIT_IN;
wire DCRPPCDSREAD_IN;
wire DCRPPCDSWRITE_IN;
wire EICC440CRITIRQ_IN;
wire EICC440EXTIRQ_IN;
wire FCMAPUCONFIRMINSTR_IN;
wire FCMAPUDONE_IN;
wire FCMAPUEXCEPTION_IN;
wire FCMAPUFPSCRFEX_IN;
wire FCMAPURESULTVALID_IN;
wire FCMAPUSLEEPNOTREADY_IN;
wire JTGC440TCK_IN;
wire JTGC440TDI_IN;
wire JTGC440TMS_IN;
wire JTGC440TRSTNEG_IN;
wire LLDMA0RSTENGINEREQ_IN;
wire LLDMA0RXEOFN_IN;
wire LLDMA0RXEOPN_IN;
wire LLDMA0RXSOFN_IN;
wire LLDMA0RXSOPN_IN;
wire LLDMA0RXSRCRDYN_IN;
wire LLDMA0TXDSTRDYN_IN;
wire LLDMA1RSTENGINEREQ_IN;
wire LLDMA1RXEOFN_IN;
wire LLDMA1RXEOPN_IN;
wire LLDMA1RXSOFN_IN;
wire LLDMA1RXSOPN_IN;
wire LLDMA1RXSRCRDYN_IN;
wire LLDMA1TXDSTRDYN_IN;
wire LLDMA2RSTENGINEREQ_IN;
wire LLDMA2RXEOFN_IN;
wire LLDMA2RXEOPN_IN;
wire LLDMA2RXSOFN_IN;
wire LLDMA2RXSOPN_IN;
wire LLDMA2RXSRCRDYN_IN;
wire LLDMA2TXDSTRDYN_IN;
wire LLDMA3RSTENGINEREQ_IN;
wire LLDMA3RXEOFN_IN;
wire LLDMA3RXEOPN_IN;
wire LLDMA3RXSOFN_IN;
wire LLDMA3RXSOPN_IN;
wire LLDMA3RXSRCRDYN_IN;
wire LLDMA3TXDSTRDYN_IN;
wire MCMIADDRREADYTOACCEPT_IN;
wire MCMIREADDATAERR_IN;
wire MCMIREADDATAVALID_IN;
wire PLBPPCMADDRACK_IN;
wire PLBPPCMMBUSY_IN;
wire PLBPPCMMIRQ_IN;
wire PLBPPCMMRDERR_IN;
wire PLBPPCMMWRERR_IN;
wire PLBPPCMRDBTERM_IN;
wire PLBPPCMRDDACK_IN;
wire PLBPPCMRDPENDREQ_IN;
wire PLBPPCMREARBITRATE_IN;
wire PLBPPCMTIMEOUT_IN;
wire PLBPPCMWRBTERM_IN;
wire PLBPPCMWRDACK_IN;
wire PLBPPCMWRPENDREQ_IN;
wire PLBPPCS0ABORT_IN;
wire PLBPPCS0BUSLOCK_IN;
wire PLBPPCS0LOCKERR_IN;
wire PLBPPCS0PAVALID_IN;
wire PLBPPCS0RDBURST_IN;
wire PLBPPCS0RDPENDREQ_IN;
wire PLBPPCS0RDPRIM_IN;
wire PLBPPCS0RNW_IN;
wire PLBPPCS0SAVALID_IN;
wire PLBPPCS0WRBURST_IN;
wire PLBPPCS0WRPENDREQ_IN;
wire PLBPPCS0WRPRIM_IN;
wire PLBPPCS1ABORT_IN;
wire PLBPPCS1BUSLOCK_IN;
wire PLBPPCS1LOCKERR_IN;
wire PLBPPCS1PAVALID_IN;
wire PLBPPCS1RDBURST_IN;
wire PLBPPCS1RDPENDREQ_IN;
wire PLBPPCS1RDPRIM_IN;
wire PLBPPCS1RNW_IN;
wire PLBPPCS1SAVALID_IN;
wire PLBPPCS1WRBURST_IN;
wire PLBPPCS1WRPENDREQ_IN;
wire PLBPPCS1WRPRIM_IN;
wire RSTC440RESETCHIP_IN;
wire RSTC440RESETCORE_IN;
wire RSTC440RESETSYSTEM_IN;
wire TIEC440ENDIANRESET_IN;
wire TRCC440TRACEDISABLE_IN;
wire TRCC440TRIGGEREVENTIN_IN;
wire [0:127] FCMAPUSTOREDATA_IN;
wire [0:127] MCMIREADDATA_IN;
wire [0:127] PLBPPCMRDDBUS_IN;
wire [0:127] PLBPPCS0WRDBUS_IN;
wire [0:127] PLBPPCS1WRDBUS_IN;
wire [0:15] PLBPPCS0BE_IN;
wire [0:15] PLBPPCS0TATTRIBUTE_IN;
wire [0:15] PLBPPCS1BE_IN;
wire [0:15] PLBPPCS1TATTRIBUTE_IN;
wire [0:1] PLBPPCMRDPENDPRI_IN;
wire [0:1] PLBPPCMREQPRI_IN;
wire [0:1] PLBPPCMSSIZE_IN;
wire [0:1] PLBPPCMWRPENDPRI_IN;
wire [0:1] PLBPPCS0MASTERID_IN;
wire [0:1] PLBPPCS0MSIZE_IN;
wire [0:1] PLBPPCS0RDPENDPRI_IN;
wire [0:1] PLBPPCS0REQPRI_IN;
wire [0:1] PLBPPCS0WRPENDPRI_IN;
wire [0:1] PLBPPCS1MASTERID_IN;
wire [0:1] PLBPPCS1MSIZE_IN;
wire [0:1] PLBPPCS1RDPENDPRI_IN;
wire [0:1] PLBPPCS1REQPRI_IN;
wire [0:1] PLBPPCS1WRPENDPRI_IN;
wire [0:1] TIEC440DCURDLDCACHEPLBPRIO_IN;
wire [0:1] TIEC440DCURDNONCACHEPLBPRIO_IN;
wire [0:1] TIEC440DCURDTOUCHPLBPRIO_IN;
wire [0:1] TIEC440DCURDURGENTPLBPRIO_IN;
wire [0:1] TIEC440DCUWRFLUSHPLBPRIO_IN;
wire [0:1] TIEC440DCUWRSTOREPLBPRIO_IN;
wire [0:1] TIEC440DCUWRURGENTPLBPRIO_IN;
wire [0:1] TIEC440ICURDFETCHPLBPRIO_IN;
wire [0:1] TIEC440ICURDSPECPLBPRIO_IN;
wire [0:1] TIEC440ICURDTOUCHPLBPRIO_IN;
wire [0:1] TIEDCRBASEADDR_IN;
wire [0:2] PLBPPCS0TYPE_IN;
wire [0:2] PLBPPCS1TYPE_IN;
wire [0:31] DCRPPCDMDBUSIN_IN;
wire [0:31] DCRPPCDSDBUSOUT_IN;
wire [0:31] FCMAPURESULT_IN;
wire [0:31] LLDMA0RXD_IN;
wire [0:31] LLDMA1RXD_IN;
wire [0:31] LLDMA2RXD_IN;
wire [0:31] LLDMA3RXD_IN;
wire [0:31] PLBPPCS0ABUS_IN;
wire [0:31] PLBPPCS1ABUS_IN;
wire [0:3] FCMAPUCR_IN;
wire [0:3] LLDMA0RXREM_IN;
wire [0:3] LLDMA1RXREM_IN;
wire [0:3] LLDMA2RXREM_IN;
wire [0:3] LLDMA3RXREM_IN;
wire [0:3] PLBPPCMRDWDADDR_IN;
wire [0:3] PLBPPCS0SIZE_IN;
wire [0:3] PLBPPCS1SIZE_IN;
wire [0:3] TIEC440ERPNRESET_IN;
wire [0:3] TIEC440USERRESET_IN;
wire [0:4] DBGC440SYSTEMSTATUS_IN;
wire [0:9] DCRPPCDSABUS_IN;
wire [28:31] PLBPPCS0UABUS_IN;
wire [28:31] PLBPPCS1UABUS_IN;
wire [28:31] TIEC440PIR_IN;
wire [28:31] TIEC440PVR_IN;



initial begin
	case (PPCS0_WIDTH_128N64)
		"FALSE" : PPCS0_WIDTH_128N64_BINARY = 1'b0;
		"TRUE" : PPCS0_WIDTH_128N64_BINARY = 1'b1;
		default : begin
			$display("Attribute Syntax Error : The Attribute PPCS0_WIDTH_128N64 on X_PPC440 instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", PPCS0_WIDTH_128N64);
			$finish;
		end
	endcase

	case (PPCS1_WIDTH_128N64)
		"FALSE" : PPCS1_WIDTH_128N64_BINARY = 1'b0;
		"TRUE" : PPCS1_WIDTH_128N64_BINARY = 1'b1;
		default : begin
			$display("Attribute Syntax Error : The Attribute PPCS1_WIDTH_128N64 on X_PPC440 instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", PPCS1_WIDTH_128N64);
			$finish;
		end
	endcase

	case (PPCDM_ASYNCMODE)
		"FALSE" : PPCDM_ASYNCMODE_BINARY = 1'b0;
		"TRUE" : PPCDM_ASYNCMODE_BINARY = 1'b1;
		default : begin
			$display("Attribute Syntax Error : The Attribute PPCDM_ASYNCMODE on X_PPC440 instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", PPCDM_ASYNCMODE);
			$finish;
		end
	endcase

	case (PPCDS_ASYNCMODE)
		"FALSE" : PPCDS_ASYNCMODE_BINARY = 1'b0;
		"TRUE" : PPCDS_ASYNCMODE_BINARY = 1'b1;
		default : begin
			$display("Attribute Syntax Error : The Attribute PPCDS_ASYNCMODE on X_PPC440 instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", PPCDS_ASYNCMODE);
			$finish;
		end
	endcase

	case (DCR_AUTOLOCK_ENABLE)
		"FALSE" : DCR_AUTOLOCK_ENABLE_BINARY = 1'b0;
		"TRUE" : DCR_AUTOLOCK_ENABLE_BINARY = 1'b1;
		default : begin
			$display("Attribute Syntax Error : The Attribute DCR_AUTOLOCK_ENABLE on X_PPC440 instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", DCR_AUTOLOCK_ENABLE);
			$finish;
		end
	endcase

	case (CLOCK_DELAY)
//		"FALSE" : CLOCK_DELAY_BINARY = 1'b0;
//		"TRUE" : CLOCK_DELAY_BINARY = 1'b1;
//		"FALSE" : CLOCK_DELAY_BINARY = 5'b00100;
		"FALSE" : CLOCK_DELAY_BINARY = 5'b10000;
		"TRUE" : CLOCK_DELAY_BINARY = 5'b00000;
		default : begin
			$display("Attribute Syntax Error : The Attribute CLOCK_DELAY on X_PPC440 instance %m is set to %s.  Legal values for this attribute are TRUE or FALSE.", CLOCK_DELAY);
			$finish;
		end
	endcase

end

buf B_DMA0LLRSTENGINEACK (DMA0LLRSTENGINEACK, DMA0LLRSTENGINEACK_OUT);
buf B_DMA0LLRXDSTRDYN (DMA0LLRXDSTRDYN, DMA0LLRXDSTRDYN_OUT);
buf B_DMA0LLTXD0 (DMA0LLTXD[0], DMA0LLTXD_OUT[0]);
buf B_DMA0LLTXD1 (DMA0LLTXD[1], DMA0LLTXD_OUT[1]);
buf B_DMA0LLTXD2 (DMA0LLTXD[2], DMA0LLTXD_OUT[2]);
buf B_DMA0LLTXD3 (DMA0LLTXD[3], DMA0LLTXD_OUT[3]);
buf B_DMA0LLTXD4 (DMA0LLTXD[4], DMA0LLTXD_OUT[4]);
buf B_DMA0LLTXD5 (DMA0LLTXD[5], DMA0LLTXD_OUT[5]);
buf B_DMA0LLTXD6 (DMA0LLTXD[6], DMA0LLTXD_OUT[6]);
buf B_DMA0LLTXD7 (DMA0LLTXD[7], DMA0LLTXD_OUT[7]);
buf B_DMA0LLTXD8 (DMA0LLTXD[8], DMA0LLTXD_OUT[8]);
buf B_DMA0LLTXD9 (DMA0LLTXD[9], DMA0LLTXD_OUT[9]);
buf B_DMA0LLTXD10 (DMA0LLTXD[10], DMA0LLTXD_OUT[10]);
buf B_DMA0LLTXD11 (DMA0LLTXD[11], DMA0LLTXD_OUT[11]);
buf B_DMA0LLTXD12 (DMA0LLTXD[12], DMA0LLTXD_OUT[12]);
buf B_DMA0LLTXD13 (DMA0LLTXD[13], DMA0LLTXD_OUT[13]);
buf B_DMA0LLTXD14 (DMA0LLTXD[14], DMA0LLTXD_OUT[14]);
buf B_DMA0LLTXD15 (DMA0LLTXD[15], DMA0LLTXD_OUT[15]);
buf B_DMA0LLTXD16 (DMA0LLTXD[16], DMA0LLTXD_OUT[16]);
buf B_DMA0LLTXD17 (DMA0LLTXD[17], DMA0LLTXD_OUT[17]);
buf B_DMA0LLTXD18 (DMA0LLTXD[18], DMA0LLTXD_OUT[18]);
buf B_DMA0LLTXD19 (DMA0LLTXD[19], DMA0LLTXD_OUT[19]);
buf B_DMA0LLTXD20 (DMA0LLTXD[20], DMA0LLTXD_OUT[20]);
buf B_DMA0LLTXD21 (DMA0LLTXD[21], DMA0LLTXD_OUT[21]);
buf B_DMA0LLTXD22 (DMA0LLTXD[22], DMA0LLTXD_OUT[22]);
buf B_DMA0LLTXD23 (DMA0LLTXD[23], DMA0LLTXD_OUT[23]);
buf B_DMA0LLTXD24 (DMA0LLTXD[24], DMA0LLTXD_OUT[24]);
buf B_DMA0LLTXD25 (DMA0LLTXD[25], DMA0LLTXD_OUT[25]);
buf B_DMA0LLTXD26 (DMA0LLTXD[26], DMA0LLTXD_OUT[26]);
buf B_DMA0LLTXD27 (DMA0LLTXD[27], DMA0LLTXD_OUT[27]);
buf B_DMA0LLTXD28 (DMA0LLTXD[28], DMA0LLTXD_OUT[28]);
buf B_DMA0LLTXD29 (DMA0LLTXD[29], DMA0LLTXD_OUT[29]);
buf B_DMA0LLTXD30 (DMA0LLTXD[30], DMA0LLTXD_OUT[30]);
buf B_DMA0LLTXD31 (DMA0LLTXD[31], DMA0LLTXD_OUT[31]);
buf B_DMA0LLTXEOFN (DMA0LLTXEOFN, DMA0LLTXEOFN_OUT);
buf B_DMA0LLTXEOPN (DMA0LLTXEOPN, DMA0LLTXEOPN_OUT);
buf B_DMA0LLTXREM0 (DMA0LLTXREM[0], DMA0LLTXREM_OUT[0]);
buf B_DMA0LLTXREM1 (DMA0LLTXREM[1], DMA0LLTXREM_OUT[1]);
buf B_DMA0LLTXREM2 (DMA0LLTXREM[2], DMA0LLTXREM_OUT[2]);
buf B_DMA0LLTXREM3 (DMA0LLTXREM[3], DMA0LLTXREM_OUT[3]);
buf B_DMA0LLTXSOFN (DMA0LLTXSOFN, DMA0LLTXSOFN_OUT);
buf B_DMA0LLTXSOPN (DMA0LLTXSOPN, DMA0LLTXSOPN_OUT);
buf B_DMA0LLTXSRCRDYN (DMA0LLTXSRCRDYN, DMA0LLTXSRCRDYN_OUT);
buf B_DMA0RXIRQ (DMA0RXIRQ, DMA0RXIRQ_OUT);
buf B_DMA0TXIRQ (DMA0TXIRQ, DMA0TXIRQ_OUT);
buf B_DMA1LLRSTENGINEACK (DMA1LLRSTENGINEACK, DMA1LLRSTENGINEACK_OUT);
buf B_DMA1LLRXDSTRDYN (DMA1LLRXDSTRDYN, DMA1LLRXDSTRDYN_OUT);
buf B_DMA1LLTXD0 (DMA1LLTXD[0], DMA1LLTXD_OUT[0]);
buf B_DMA1LLTXD1 (DMA1LLTXD[1], DMA1LLTXD_OUT[1]);
buf B_DMA1LLTXD2 (DMA1LLTXD[2], DMA1LLTXD_OUT[2]);
buf B_DMA1LLTXD3 (DMA1LLTXD[3], DMA1LLTXD_OUT[3]);
buf B_DMA1LLTXD4 (DMA1LLTXD[4], DMA1LLTXD_OUT[4]);
buf B_DMA1LLTXD5 (DMA1LLTXD[5], DMA1LLTXD_OUT[5]);
buf B_DMA1LLTXD6 (DMA1LLTXD[6], DMA1LLTXD_OUT[6]);
buf B_DMA1LLTXD7 (DMA1LLTXD[7], DMA1LLTXD_OUT[7]);
buf B_DMA1LLTXD8 (DMA1LLTXD[8], DMA1LLTXD_OUT[8]);
buf B_DMA1LLTXD9 (DMA1LLTXD[9], DMA1LLTXD_OUT[9]);
buf B_DMA1LLTXD10 (DMA1LLTXD[10], DMA1LLTXD_OUT[10]);
buf B_DMA1LLTXD11 (DMA1LLTXD[11], DMA1LLTXD_OUT[11]);
buf B_DMA1LLTXD12 (DMA1LLTXD[12], DMA1LLTXD_OUT[12]);
buf B_DMA1LLTXD13 (DMA1LLTXD[13], DMA1LLTXD_OUT[13]);
buf B_DMA1LLTXD14 (DMA1LLTXD[14], DMA1LLTXD_OUT[14]);
buf B_DMA1LLTXD15 (DMA1LLTXD[15], DMA1LLTXD_OUT[15]);
buf B_DMA1LLTXD16 (DMA1LLTXD[16], DMA1LLTXD_OUT[16]);
buf B_DMA1LLTXD17 (DMA1LLTXD[17], DMA1LLTXD_OUT[17]);
buf B_DMA1LLTXD18 (DMA1LLTXD[18], DMA1LLTXD_OUT[18]);
buf B_DMA1LLTXD19 (DMA1LLTXD[19], DMA1LLTXD_OUT[19]);
buf B_DMA1LLTXD20 (DMA1LLTXD[20], DMA1LLTXD_OUT[20]);
buf B_DMA1LLTXD21 (DMA1LLTXD[21], DMA1LLTXD_OUT[21]);
buf B_DMA1LLTXD22 (DMA1LLTXD[22], DMA1LLTXD_OUT[22]);
buf B_DMA1LLTXD23 (DMA1LLTXD[23], DMA1LLTXD_OUT[23]);
buf B_DMA1LLTXD24 (DMA1LLTXD[24], DMA1LLTXD_OUT[24]);
buf B_DMA1LLTXD25 (DMA1LLTXD[25], DMA1LLTXD_OUT[25]);
buf B_DMA1LLTXD26 (DMA1LLTXD[26], DMA1LLTXD_OUT[26]);
buf B_DMA1LLTXD27 (DMA1LLTXD[27], DMA1LLTXD_OUT[27]);
buf B_DMA1LLTXD28 (DMA1LLTXD[28], DMA1LLTXD_OUT[28]);
buf B_DMA1LLTXD29 (DMA1LLTXD[29], DMA1LLTXD_OUT[29]);
buf B_DMA1LLTXD30 (DMA1LLTXD[30], DMA1LLTXD_OUT[30]);
buf B_DMA1LLTXD31 (DMA1LLTXD[31], DMA1LLTXD_OUT[31]);
buf B_DMA1LLTXEOFN (DMA1LLTXEOFN, DMA1LLTXEOFN_OUT);
buf B_DMA1LLTXEOPN (DMA1LLTXEOPN, DMA1LLTXEOPN_OUT);
buf B_DMA1LLTXREM0 (DMA1LLTXREM[0], DMA1LLTXREM_OUT[0]);
buf B_DMA1LLTXREM1 (DMA1LLTXREM[1], DMA1LLTXREM_OUT[1]);
buf B_DMA1LLTXREM2 (DMA1LLTXREM[2], DMA1LLTXREM_OUT[2]);
buf B_DMA1LLTXREM3 (DMA1LLTXREM[3], DMA1LLTXREM_OUT[3]);
buf B_DMA1LLTXSOFN (DMA1LLTXSOFN, DMA1LLTXSOFN_OUT);
buf B_DMA1LLTXSOPN (DMA1LLTXSOPN, DMA1LLTXSOPN_OUT);
buf B_DMA1LLTXSRCRDYN (DMA1LLTXSRCRDYN, DMA1LLTXSRCRDYN_OUT);
buf B_DMA1RXIRQ (DMA1RXIRQ, DMA1RXIRQ_OUT);
buf B_DMA1TXIRQ (DMA1TXIRQ, DMA1TXIRQ_OUT);
buf B_DMA2LLRSTENGINEACK (DMA2LLRSTENGINEACK, DMA2LLRSTENGINEACK_OUT);
buf B_DMA2LLRXDSTRDYN (DMA2LLRXDSTRDYN, DMA2LLRXDSTRDYN_OUT);
buf B_DMA2LLTXD0 (DMA2LLTXD[0], DMA2LLTXD_OUT[0]);
buf B_DMA2LLTXD1 (DMA2LLTXD[1], DMA2LLTXD_OUT[1]);
buf B_DMA2LLTXD2 (DMA2LLTXD[2], DMA2LLTXD_OUT[2]);
buf B_DMA2LLTXD3 (DMA2LLTXD[3], DMA2LLTXD_OUT[3]);
buf B_DMA2LLTXD4 (DMA2LLTXD[4], DMA2LLTXD_OUT[4]);
buf B_DMA2LLTXD5 (DMA2LLTXD[5], DMA2LLTXD_OUT[5]);
buf B_DMA2LLTXD6 (DMA2LLTXD[6], DMA2LLTXD_OUT[6]);
buf B_DMA2LLTXD7 (DMA2LLTXD[7], DMA2LLTXD_OUT[7]);
buf B_DMA2LLTXD8 (DMA2LLTXD[8], DMA2LLTXD_OUT[8]);
buf B_DMA2LLTXD9 (DMA2LLTXD[9], DMA2LLTXD_OUT[9]);
buf B_DMA2LLTXD10 (DMA2LLTXD[10], DMA2LLTXD_OUT[10]);
buf B_DMA2LLTXD11 (DMA2LLTXD[11], DMA2LLTXD_OUT[11]);
buf B_DMA2LLTXD12 (DMA2LLTXD[12], DMA2LLTXD_OUT[12]);
buf B_DMA2LLTXD13 (DMA2LLTXD[13], DMA2LLTXD_OUT[13]);
buf B_DMA2LLTXD14 (DMA2LLTXD[14], DMA2LLTXD_OUT[14]);
buf B_DMA2LLTXD15 (DMA2LLTXD[15], DMA2LLTXD_OUT[15]);
buf B_DMA2LLTXD16 (DMA2LLTXD[16], DMA2LLTXD_OUT[16]);
buf B_DMA2LLTXD17 (DMA2LLTXD[17], DMA2LLTXD_OUT[17]);
buf B_DMA2LLTXD18 (DMA2LLTXD[18], DMA2LLTXD_OUT[18]);
buf B_DMA2LLTXD19 (DMA2LLTXD[19], DMA2LLTXD_OUT[19]);
buf B_DMA2LLTXD20 (DMA2LLTXD[20], DMA2LLTXD_OUT[20]);
buf B_DMA2LLTXD21 (DMA2LLTXD[21], DMA2LLTXD_OUT[21]);
buf B_DMA2LLTXD22 (DMA2LLTXD[22], DMA2LLTXD_OUT[22]);
buf B_DMA2LLTXD23 (DMA2LLTXD[23], DMA2LLTXD_OUT[23]);
buf B_DMA2LLTXD24 (DMA2LLTXD[24], DMA2LLTXD_OUT[24]);
buf B_DMA2LLTXD25 (DMA2LLTXD[25], DMA2LLTXD_OUT[25]);
buf B_DMA2LLTXD26 (DMA2LLTXD[26], DMA2LLTXD_OUT[26]);
buf B_DMA2LLTXD27 (DMA2LLTXD[27], DMA2LLTXD_OUT[27]);
buf B_DMA2LLTXD28 (DMA2LLTXD[28], DMA2LLTXD_OUT[28]);
buf B_DMA2LLTXD29 (DMA2LLTXD[29], DMA2LLTXD_OUT[29]);
buf B_DMA2LLTXD30 (DMA2LLTXD[30], DMA2LLTXD_OUT[30]);
buf B_DMA2LLTXD31 (DMA2LLTXD[31], DMA2LLTXD_OUT[31]);
buf B_DMA2LLTXEOFN (DMA2LLTXEOFN, DMA2LLTXEOFN_OUT);
buf B_DMA2LLTXEOPN (DMA2LLTXEOPN, DMA2LLTXEOPN_OUT);
buf B_DMA2LLTXREM0 (DMA2LLTXREM[0], DMA2LLTXREM_OUT[0]);
buf B_DMA2LLTXREM1 (DMA2LLTXREM[1], DMA2LLTXREM_OUT[1]);
buf B_DMA2LLTXREM2 (DMA2LLTXREM[2], DMA2LLTXREM_OUT[2]);
buf B_DMA2LLTXREM3 (DMA2LLTXREM[3], DMA2LLTXREM_OUT[3]);
buf B_DMA2LLTXSOFN (DMA2LLTXSOFN, DMA2LLTXSOFN_OUT);
buf B_DMA2LLTXSOPN (DMA2LLTXSOPN, DMA2LLTXSOPN_OUT);
buf B_DMA2LLTXSRCRDYN (DMA2LLTXSRCRDYN, DMA2LLTXSRCRDYN_OUT);
buf B_DMA2RXIRQ (DMA2RXIRQ, DMA2RXIRQ_OUT);
buf B_DMA2TXIRQ (DMA2TXIRQ, DMA2TXIRQ_OUT);
buf B_DMA3LLRSTENGINEACK (DMA3LLRSTENGINEACK, DMA3LLRSTENGINEACK_OUT);
buf B_DMA3LLRXDSTRDYN (DMA3LLRXDSTRDYN, DMA3LLRXDSTRDYN_OUT);
buf B_DMA3LLTXD0 (DMA3LLTXD[0], DMA3LLTXD_OUT[0]);
buf B_DMA3LLTXD1 (DMA3LLTXD[1], DMA3LLTXD_OUT[1]);
buf B_DMA3LLTXD2 (DMA3LLTXD[2], DMA3LLTXD_OUT[2]);
buf B_DMA3LLTXD3 (DMA3LLTXD[3], DMA3LLTXD_OUT[3]);
buf B_DMA3LLTXD4 (DMA3LLTXD[4], DMA3LLTXD_OUT[4]);
buf B_DMA3LLTXD5 (DMA3LLTXD[5], DMA3LLTXD_OUT[5]);
buf B_DMA3LLTXD6 (DMA3LLTXD[6], DMA3LLTXD_OUT[6]);
buf B_DMA3LLTXD7 (DMA3LLTXD[7], DMA3LLTXD_OUT[7]);
buf B_DMA3LLTXD8 (DMA3LLTXD[8], DMA3LLTXD_OUT[8]);
buf B_DMA3LLTXD9 (DMA3LLTXD[9], DMA3LLTXD_OUT[9]);
buf B_DMA3LLTXD10 (DMA3LLTXD[10], DMA3LLTXD_OUT[10]);
buf B_DMA3LLTXD11 (DMA3LLTXD[11], DMA3LLTXD_OUT[11]);
buf B_DMA3LLTXD12 (DMA3LLTXD[12], DMA3LLTXD_OUT[12]);
buf B_DMA3LLTXD13 (DMA3LLTXD[13], DMA3LLTXD_OUT[13]);
buf B_DMA3LLTXD14 (DMA3LLTXD[14], DMA3LLTXD_OUT[14]);
buf B_DMA3LLTXD15 (DMA3LLTXD[15], DMA3LLTXD_OUT[15]);
buf B_DMA3LLTXD16 (DMA3LLTXD[16], DMA3LLTXD_OUT[16]);
buf B_DMA3LLTXD17 (DMA3LLTXD[17], DMA3LLTXD_OUT[17]);
buf B_DMA3LLTXD18 (DMA3LLTXD[18], DMA3LLTXD_OUT[18]);
buf B_DMA3LLTXD19 (DMA3LLTXD[19], DMA3LLTXD_OUT[19]);
buf B_DMA3LLTXD20 (DMA3LLTXD[20], DMA3LLTXD_OUT[20]);
buf B_DMA3LLTXD21 (DMA3LLTXD[21], DMA3LLTXD_OUT[21]);
buf B_DMA3LLTXD22 (DMA3LLTXD[22], DMA3LLTXD_OUT[22]);
buf B_DMA3LLTXD23 (DMA3LLTXD[23], DMA3LLTXD_OUT[23]);
buf B_DMA3LLTXD24 (DMA3LLTXD[24], DMA3LLTXD_OUT[24]);
buf B_DMA3LLTXD25 (DMA3LLTXD[25], DMA3LLTXD_OUT[25]);
buf B_DMA3LLTXD26 (DMA3LLTXD[26], DMA3LLTXD_OUT[26]);
buf B_DMA3LLTXD27 (DMA3LLTXD[27], DMA3LLTXD_OUT[27]);
buf B_DMA3LLTXD28 (DMA3LLTXD[28], DMA3LLTXD_OUT[28]);
buf B_DMA3LLTXD29 (DMA3LLTXD[29], DMA3LLTXD_OUT[29]);
buf B_DMA3LLTXD30 (DMA3LLTXD[30], DMA3LLTXD_OUT[30]);
buf B_DMA3LLTXD31 (DMA3LLTXD[31], DMA3LLTXD_OUT[31]);
buf B_DMA3LLTXEOFN (DMA3LLTXEOFN, DMA3LLTXEOFN_OUT);
buf B_DMA3LLTXEOPN (DMA3LLTXEOPN, DMA3LLTXEOPN_OUT);
buf B_DMA3LLTXREM0 (DMA3LLTXREM[0], DMA3LLTXREM_OUT[0]);
buf B_DMA3LLTXREM1 (DMA3LLTXREM[1], DMA3LLTXREM_OUT[1]);
buf B_DMA3LLTXREM2 (DMA3LLTXREM[2], DMA3LLTXREM_OUT[2]);
buf B_DMA3LLTXREM3 (DMA3LLTXREM[3], DMA3LLTXREM_OUT[3]);
buf B_DMA3LLTXSOFN (DMA3LLTXSOFN, DMA3LLTXSOFN_OUT);
buf B_DMA3LLTXSOPN (DMA3LLTXSOPN, DMA3LLTXSOPN_OUT);
buf B_DMA3LLTXSRCRDYN (DMA3LLTXSRCRDYN, DMA3LLTXSRCRDYN_OUT);
buf B_DMA3RXIRQ (DMA3RXIRQ, DMA3RXIRQ_OUT);
buf B_DMA3TXIRQ (DMA3TXIRQ, DMA3TXIRQ_OUT);
buf B_PPCDMDCRABUS0 (PPCDMDCRABUS[0], PPCDMDCRABUS_OUT[0]);
buf B_PPCDMDCRABUS1 (PPCDMDCRABUS[1], PPCDMDCRABUS_OUT[1]);
buf B_PPCDMDCRABUS2 (PPCDMDCRABUS[2], PPCDMDCRABUS_OUT[2]);
buf B_PPCDMDCRABUS3 (PPCDMDCRABUS[3], PPCDMDCRABUS_OUT[3]);
buf B_PPCDMDCRABUS4 (PPCDMDCRABUS[4], PPCDMDCRABUS_OUT[4]);
buf B_PPCDMDCRABUS5 (PPCDMDCRABUS[5], PPCDMDCRABUS_OUT[5]);
buf B_PPCDMDCRABUS6 (PPCDMDCRABUS[6], PPCDMDCRABUS_OUT[6]);
buf B_PPCDMDCRABUS7 (PPCDMDCRABUS[7], PPCDMDCRABUS_OUT[7]);
buf B_PPCDMDCRABUS8 (PPCDMDCRABUS[8], PPCDMDCRABUS_OUT[8]);
buf B_PPCDMDCRABUS9 (PPCDMDCRABUS[9], PPCDMDCRABUS_OUT[9]);
buf B_PPCDMDCRDBUSOUT0 (PPCDMDCRDBUSOUT[0], PPCDMDCRDBUSOUT_OUT[0]);
buf B_PPCDMDCRDBUSOUT1 (PPCDMDCRDBUSOUT[1], PPCDMDCRDBUSOUT_OUT[1]);
buf B_PPCDMDCRDBUSOUT2 (PPCDMDCRDBUSOUT[2], PPCDMDCRDBUSOUT_OUT[2]);
buf B_PPCDMDCRDBUSOUT3 (PPCDMDCRDBUSOUT[3], PPCDMDCRDBUSOUT_OUT[3]);
buf B_PPCDMDCRDBUSOUT4 (PPCDMDCRDBUSOUT[4], PPCDMDCRDBUSOUT_OUT[4]);
buf B_PPCDMDCRDBUSOUT5 (PPCDMDCRDBUSOUT[5], PPCDMDCRDBUSOUT_OUT[5]);
buf B_PPCDMDCRDBUSOUT6 (PPCDMDCRDBUSOUT[6], PPCDMDCRDBUSOUT_OUT[6]);
buf B_PPCDMDCRDBUSOUT7 (PPCDMDCRDBUSOUT[7], PPCDMDCRDBUSOUT_OUT[7]);
buf B_PPCDMDCRDBUSOUT8 (PPCDMDCRDBUSOUT[8], PPCDMDCRDBUSOUT_OUT[8]);
buf B_PPCDMDCRDBUSOUT9 (PPCDMDCRDBUSOUT[9], PPCDMDCRDBUSOUT_OUT[9]);
buf B_PPCDMDCRDBUSOUT10 (PPCDMDCRDBUSOUT[10], PPCDMDCRDBUSOUT_OUT[10]);
buf B_PPCDMDCRDBUSOUT11 (PPCDMDCRDBUSOUT[11], PPCDMDCRDBUSOUT_OUT[11]);
buf B_PPCDMDCRDBUSOUT12 (PPCDMDCRDBUSOUT[12], PPCDMDCRDBUSOUT_OUT[12]);
buf B_PPCDMDCRDBUSOUT13 (PPCDMDCRDBUSOUT[13], PPCDMDCRDBUSOUT_OUT[13]);
buf B_PPCDMDCRDBUSOUT14 (PPCDMDCRDBUSOUT[14], PPCDMDCRDBUSOUT_OUT[14]);
buf B_PPCDMDCRDBUSOUT15 (PPCDMDCRDBUSOUT[15], PPCDMDCRDBUSOUT_OUT[15]);
buf B_PPCDMDCRDBUSOUT16 (PPCDMDCRDBUSOUT[16], PPCDMDCRDBUSOUT_OUT[16]);
buf B_PPCDMDCRDBUSOUT17 (PPCDMDCRDBUSOUT[17], PPCDMDCRDBUSOUT_OUT[17]);
buf B_PPCDMDCRDBUSOUT18 (PPCDMDCRDBUSOUT[18], PPCDMDCRDBUSOUT_OUT[18]);
buf B_PPCDMDCRDBUSOUT19 (PPCDMDCRDBUSOUT[19], PPCDMDCRDBUSOUT_OUT[19]);
buf B_PPCDMDCRDBUSOUT20 (PPCDMDCRDBUSOUT[20], PPCDMDCRDBUSOUT_OUT[20]);
buf B_PPCDMDCRDBUSOUT21 (PPCDMDCRDBUSOUT[21], PPCDMDCRDBUSOUT_OUT[21]);
buf B_PPCDMDCRDBUSOUT22 (PPCDMDCRDBUSOUT[22], PPCDMDCRDBUSOUT_OUT[22]);
buf B_PPCDMDCRDBUSOUT23 (PPCDMDCRDBUSOUT[23], PPCDMDCRDBUSOUT_OUT[23]);
buf B_PPCDMDCRDBUSOUT24 (PPCDMDCRDBUSOUT[24], PPCDMDCRDBUSOUT_OUT[24]);
buf B_PPCDMDCRDBUSOUT25 (PPCDMDCRDBUSOUT[25], PPCDMDCRDBUSOUT_OUT[25]);
buf B_PPCDMDCRDBUSOUT26 (PPCDMDCRDBUSOUT[26], PPCDMDCRDBUSOUT_OUT[26]);
buf B_PPCDMDCRDBUSOUT27 (PPCDMDCRDBUSOUT[27], PPCDMDCRDBUSOUT_OUT[27]);
buf B_PPCDMDCRDBUSOUT28 (PPCDMDCRDBUSOUT[28], PPCDMDCRDBUSOUT_OUT[28]);
buf B_PPCDMDCRDBUSOUT29 (PPCDMDCRDBUSOUT[29], PPCDMDCRDBUSOUT_OUT[29]);
buf B_PPCDMDCRDBUSOUT30 (PPCDMDCRDBUSOUT[30], PPCDMDCRDBUSOUT_OUT[30]);
buf B_PPCDMDCRDBUSOUT31 (PPCDMDCRDBUSOUT[31], PPCDMDCRDBUSOUT_OUT[31]);
buf B_PPCDMDCRREAD (PPCDMDCRREAD, PPCDMDCRREAD_OUT);
buf B_PPCDMDCRUABUS20 (PPCDMDCRUABUS[20], PPCDMDCRUABUS_OUT[20]);
buf B_PPCDMDCRUABUS21 (PPCDMDCRUABUS[21], PPCDMDCRUABUS_OUT[21]);
buf B_PPCDMDCRWRITE (PPCDMDCRWRITE, PPCDMDCRWRITE_OUT);
buf B_PPCMPLBABORT (PPCMPLBABORT, PPCMPLBABORT_OUT);
buf B_PPCMPLBABUS0 (PPCMPLBABUS[0], PPCMPLBABUS_OUT[0]);
buf B_PPCMPLBABUS1 (PPCMPLBABUS[1], PPCMPLBABUS_OUT[1]);
buf B_PPCMPLBABUS2 (PPCMPLBABUS[2], PPCMPLBABUS_OUT[2]);
buf B_PPCMPLBABUS3 (PPCMPLBABUS[3], PPCMPLBABUS_OUT[3]);
buf B_PPCMPLBABUS4 (PPCMPLBABUS[4], PPCMPLBABUS_OUT[4]);
buf B_PPCMPLBABUS5 (PPCMPLBABUS[5], PPCMPLBABUS_OUT[5]);
buf B_PPCMPLBABUS6 (PPCMPLBABUS[6], PPCMPLBABUS_OUT[6]);
buf B_PPCMPLBABUS7 (PPCMPLBABUS[7], PPCMPLBABUS_OUT[7]);
buf B_PPCMPLBABUS8 (PPCMPLBABUS[8], PPCMPLBABUS_OUT[8]);
buf B_PPCMPLBABUS9 (PPCMPLBABUS[9], PPCMPLBABUS_OUT[9]);
buf B_PPCMPLBABUS10 (PPCMPLBABUS[10], PPCMPLBABUS_OUT[10]);
buf B_PPCMPLBABUS11 (PPCMPLBABUS[11], PPCMPLBABUS_OUT[11]);
buf B_PPCMPLBABUS12 (PPCMPLBABUS[12], PPCMPLBABUS_OUT[12]);
buf B_PPCMPLBABUS13 (PPCMPLBABUS[13], PPCMPLBABUS_OUT[13]);
buf B_PPCMPLBABUS14 (PPCMPLBABUS[14], PPCMPLBABUS_OUT[14]);
buf B_PPCMPLBABUS15 (PPCMPLBABUS[15], PPCMPLBABUS_OUT[15]);
buf B_PPCMPLBABUS16 (PPCMPLBABUS[16], PPCMPLBABUS_OUT[16]);
buf B_PPCMPLBABUS17 (PPCMPLBABUS[17], PPCMPLBABUS_OUT[17]);
buf B_PPCMPLBABUS18 (PPCMPLBABUS[18], PPCMPLBABUS_OUT[18]);
buf B_PPCMPLBABUS19 (PPCMPLBABUS[19], PPCMPLBABUS_OUT[19]);
buf B_PPCMPLBABUS20 (PPCMPLBABUS[20], PPCMPLBABUS_OUT[20]);
buf B_PPCMPLBABUS21 (PPCMPLBABUS[21], PPCMPLBABUS_OUT[21]);
buf B_PPCMPLBABUS22 (PPCMPLBABUS[22], PPCMPLBABUS_OUT[22]);
buf B_PPCMPLBABUS23 (PPCMPLBABUS[23], PPCMPLBABUS_OUT[23]);
buf B_PPCMPLBABUS24 (PPCMPLBABUS[24], PPCMPLBABUS_OUT[24]);
buf B_PPCMPLBABUS25 (PPCMPLBABUS[25], PPCMPLBABUS_OUT[25]);
buf B_PPCMPLBABUS26 (PPCMPLBABUS[26], PPCMPLBABUS_OUT[26]);
buf B_PPCMPLBABUS27 (PPCMPLBABUS[27], PPCMPLBABUS_OUT[27]);
buf B_PPCMPLBABUS28 (PPCMPLBABUS[28], PPCMPLBABUS_OUT[28]);
buf B_PPCMPLBABUS29 (PPCMPLBABUS[29], PPCMPLBABUS_OUT[29]);
buf B_PPCMPLBABUS30 (PPCMPLBABUS[30], PPCMPLBABUS_OUT[30]);
buf B_PPCMPLBABUS31 (PPCMPLBABUS[31], PPCMPLBABUS_OUT[31]);
buf B_PPCMPLBBE0 (PPCMPLBBE[0], PPCMPLBBE_OUT[0]);
buf B_PPCMPLBBE1 (PPCMPLBBE[1], PPCMPLBBE_OUT[1]);
buf B_PPCMPLBBE2 (PPCMPLBBE[2], PPCMPLBBE_OUT[2]);
buf B_PPCMPLBBE3 (PPCMPLBBE[3], PPCMPLBBE_OUT[3]);
buf B_PPCMPLBBE4 (PPCMPLBBE[4], PPCMPLBBE_OUT[4]);
buf B_PPCMPLBBE5 (PPCMPLBBE[5], PPCMPLBBE_OUT[5]);
buf B_PPCMPLBBE6 (PPCMPLBBE[6], PPCMPLBBE_OUT[6]);
buf B_PPCMPLBBE7 (PPCMPLBBE[7], PPCMPLBBE_OUT[7]);
buf B_PPCMPLBBE8 (PPCMPLBBE[8], PPCMPLBBE_OUT[8]);
buf B_PPCMPLBBE9 (PPCMPLBBE[9], PPCMPLBBE_OUT[9]);
buf B_PPCMPLBBE10 (PPCMPLBBE[10], PPCMPLBBE_OUT[10]);
buf B_PPCMPLBBE11 (PPCMPLBBE[11], PPCMPLBBE_OUT[11]);
buf B_PPCMPLBBE12 (PPCMPLBBE[12], PPCMPLBBE_OUT[12]);
buf B_PPCMPLBBE13 (PPCMPLBBE[13], PPCMPLBBE_OUT[13]);
buf B_PPCMPLBBE14 (PPCMPLBBE[14], PPCMPLBBE_OUT[14]);
buf B_PPCMPLBBE15 (PPCMPLBBE[15], PPCMPLBBE_OUT[15]);
buf B_PPCMPLBBUSLOCK (PPCMPLBBUSLOCK, PPCMPLBBUSLOCK_OUT);
buf B_PPCMPLBLOCKERR (PPCMPLBLOCKERR, PPCMPLBLOCKERR_OUT);
buf B_PPCMPLBPRIORITY0 (PPCMPLBPRIORITY[0], PPCMPLBPRIORITY_OUT[0]);
buf B_PPCMPLBPRIORITY1 (PPCMPLBPRIORITY[1], PPCMPLBPRIORITY_OUT[1]);
buf B_PPCMPLBRDBURST (PPCMPLBRDBURST, PPCMPLBRDBURST_OUT);
buf B_PPCMPLBREQUEST (PPCMPLBREQUEST, PPCMPLBREQUEST_OUT);
buf B_PPCMPLBRNW (PPCMPLBRNW, PPCMPLBRNW_OUT);
buf B_PPCMPLBSIZE0 (PPCMPLBSIZE[0], PPCMPLBSIZE_OUT[0]);
buf B_PPCMPLBSIZE1 (PPCMPLBSIZE[1], PPCMPLBSIZE_OUT[1]);
buf B_PPCMPLBSIZE2 (PPCMPLBSIZE[2], PPCMPLBSIZE_OUT[2]);
buf B_PPCMPLBSIZE3 (PPCMPLBSIZE[3], PPCMPLBSIZE_OUT[3]);
buf B_PPCMPLBTATTRIBUTE0 (PPCMPLBTATTRIBUTE[0], PPCMPLBTATTRIBUTE_OUT[0]);
buf B_PPCMPLBTATTRIBUTE1 (PPCMPLBTATTRIBUTE[1], PPCMPLBTATTRIBUTE_OUT[1]);
buf B_PPCMPLBTATTRIBUTE2 (PPCMPLBTATTRIBUTE[2], PPCMPLBTATTRIBUTE_OUT[2]);
buf B_PPCMPLBTATTRIBUTE3 (PPCMPLBTATTRIBUTE[3], PPCMPLBTATTRIBUTE_OUT[3]);
buf B_PPCMPLBTATTRIBUTE4 (PPCMPLBTATTRIBUTE[4], PPCMPLBTATTRIBUTE_OUT[4]);
buf B_PPCMPLBTATTRIBUTE5 (PPCMPLBTATTRIBUTE[5], PPCMPLBTATTRIBUTE_OUT[5]);
buf B_PPCMPLBTATTRIBUTE6 (PPCMPLBTATTRIBUTE[6], PPCMPLBTATTRIBUTE_OUT[6]);
buf B_PPCMPLBTATTRIBUTE7 (PPCMPLBTATTRIBUTE[7], PPCMPLBTATTRIBUTE_OUT[7]);
buf B_PPCMPLBTATTRIBUTE8 (PPCMPLBTATTRIBUTE[8], PPCMPLBTATTRIBUTE_OUT[8]);
buf B_PPCMPLBTATTRIBUTE9 (PPCMPLBTATTRIBUTE[9], PPCMPLBTATTRIBUTE_OUT[9]);
buf B_PPCMPLBTATTRIBUTE10 (PPCMPLBTATTRIBUTE[10], PPCMPLBTATTRIBUTE_OUT[10]);
buf B_PPCMPLBTATTRIBUTE11 (PPCMPLBTATTRIBUTE[11], PPCMPLBTATTRIBUTE_OUT[11]);
buf B_PPCMPLBTATTRIBUTE12 (PPCMPLBTATTRIBUTE[12], PPCMPLBTATTRIBUTE_OUT[12]);
buf B_PPCMPLBTATTRIBUTE13 (PPCMPLBTATTRIBUTE[13], PPCMPLBTATTRIBUTE_OUT[13]);
buf B_PPCMPLBTATTRIBUTE14 (PPCMPLBTATTRIBUTE[14], PPCMPLBTATTRIBUTE_OUT[14]);
buf B_PPCMPLBTATTRIBUTE15 (PPCMPLBTATTRIBUTE[15], PPCMPLBTATTRIBUTE_OUT[15]);
buf B_PPCMPLBTYPE0 (PPCMPLBTYPE[0], PPCMPLBTYPE_OUT[0]);
buf B_PPCMPLBTYPE1 (PPCMPLBTYPE[1], PPCMPLBTYPE_OUT[1]);
buf B_PPCMPLBTYPE2 (PPCMPLBTYPE[2], PPCMPLBTYPE_OUT[2]);
buf B_PPCMPLBUABUS28 (PPCMPLBUABUS[28], PPCMPLBUABUS_OUT[28]);
buf B_PPCMPLBUABUS29 (PPCMPLBUABUS[29], PPCMPLBUABUS_OUT[29]);
buf B_PPCMPLBUABUS30 (PPCMPLBUABUS[30], PPCMPLBUABUS_OUT[30]);
buf B_PPCMPLBUABUS31 (PPCMPLBUABUS[31], PPCMPLBUABUS_OUT[31]);
buf B_PPCMPLBWRBURST (PPCMPLBWRBURST, PPCMPLBWRBURST_OUT);
buf B_PPCMPLBWRDBUS0 (PPCMPLBWRDBUS[0], PPCMPLBWRDBUS_OUT[0]);
buf B_PPCMPLBWRDBUS1 (PPCMPLBWRDBUS[1], PPCMPLBWRDBUS_OUT[1]);
buf B_PPCMPLBWRDBUS2 (PPCMPLBWRDBUS[2], PPCMPLBWRDBUS_OUT[2]);
buf B_PPCMPLBWRDBUS3 (PPCMPLBWRDBUS[3], PPCMPLBWRDBUS_OUT[3]);
buf B_PPCMPLBWRDBUS4 (PPCMPLBWRDBUS[4], PPCMPLBWRDBUS_OUT[4]);
buf B_PPCMPLBWRDBUS5 (PPCMPLBWRDBUS[5], PPCMPLBWRDBUS_OUT[5]);
buf B_PPCMPLBWRDBUS6 (PPCMPLBWRDBUS[6], PPCMPLBWRDBUS_OUT[6]);
buf B_PPCMPLBWRDBUS7 (PPCMPLBWRDBUS[7], PPCMPLBWRDBUS_OUT[7]);
buf B_PPCMPLBWRDBUS8 (PPCMPLBWRDBUS[8], PPCMPLBWRDBUS_OUT[8]);
buf B_PPCMPLBWRDBUS9 (PPCMPLBWRDBUS[9], PPCMPLBWRDBUS_OUT[9]);
buf B_PPCMPLBWRDBUS10 (PPCMPLBWRDBUS[10], PPCMPLBWRDBUS_OUT[10]);
buf B_PPCMPLBWRDBUS11 (PPCMPLBWRDBUS[11], PPCMPLBWRDBUS_OUT[11]);
buf B_PPCMPLBWRDBUS12 (PPCMPLBWRDBUS[12], PPCMPLBWRDBUS_OUT[12]);
buf B_PPCMPLBWRDBUS13 (PPCMPLBWRDBUS[13], PPCMPLBWRDBUS_OUT[13]);
buf B_PPCMPLBWRDBUS14 (PPCMPLBWRDBUS[14], PPCMPLBWRDBUS_OUT[14]);
buf B_PPCMPLBWRDBUS15 (PPCMPLBWRDBUS[15], PPCMPLBWRDBUS_OUT[15]);
buf B_PPCMPLBWRDBUS16 (PPCMPLBWRDBUS[16], PPCMPLBWRDBUS_OUT[16]);
buf B_PPCMPLBWRDBUS17 (PPCMPLBWRDBUS[17], PPCMPLBWRDBUS_OUT[17]);
buf B_PPCMPLBWRDBUS18 (PPCMPLBWRDBUS[18], PPCMPLBWRDBUS_OUT[18]);
buf B_PPCMPLBWRDBUS19 (PPCMPLBWRDBUS[19], PPCMPLBWRDBUS_OUT[19]);
buf B_PPCMPLBWRDBUS20 (PPCMPLBWRDBUS[20], PPCMPLBWRDBUS_OUT[20]);
buf B_PPCMPLBWRDBUS21 (PPCMPLBWRDBUS[21], PPCMPLBWRDBUS_OUT[21]);
buf B_PPCMPLBWRDBUS22 (PPCMPLBWRDBUS[22], PPCMPLBWRDBUS_OUT[22]);
buf B_PPCMPLBWRDBUS23 (PPCMPLBWRDBUS[23], PPCMPLBWRDBUS_OUT[23]);
buf B_PPCMPLBWRDBUS24 (PPCMPLBWRDBUS[24], PPCMPLBWRDBUS_OUT[24]);
buf B_PPCMPLBWRDBUS25 (PPCMPLBWRDBUS[25], PPCMPLBWRDBUS_OUT[25]);
buf B_PPCMPLBWRDBUS26 (PPCMPLBWRDBUS[26], PPCMPLBWRDBUS_OUT[26]);
buf B_PPCMPLBWRDBUS27 (PPCMPLBWRDBUS[27], PPCMPLBWRDBUS_OUT[27]);
buf B_PPCMPLBWRDBUS28 (PPCMPLBWRDBUS[28], PPCMPLBWRDBUS_OUT[28]);
buf B_PPCMPLBWRDBUS29 (PPCMPLBWRDBUS[29], PPCMPLBWRDBUS_OUT[29]);
buf B_PPCMPLBWRDBUS30 (PPCMPLBWRDBUS[30], PPCMPLBWRDBUS_OUT[30]);
buf B_PPCMPLBWRDBUS31 (PPCMPLBWRDBUS[31], PPCMPLBWRDBUS_OUT[31]);
buf B_PPCMPLBWRDBUS32 (PPCMPLBWRDBUS[32], PPCMPLBWRDBUS_OUT[32]);
buf B_PPCMPLBWRDBUS33 (PPCMPLBWRDBUS[33], PPCMPLBWRDBUS_OUT[33]);
buf B_PPCMPLBWRDBUS34 (PPCMPLBWRDBUS[34], PPCMPLBWRDBUS_OUT[34]);
buf B_PPCMPLBWRDBUS35 (PPCMPLBWRDBUS[35], PPCMPLBWRDBUS_OUT[35]);
buf B_PPCMPLBWRDBUS36 (PPCMPLBWRDBUS[36], PPCMPLBWRDBUS_OUT[36]);
buf B_PPCMPLBWRDBUS37 (PPCMPLBWRDBUS[37], PPCMPLBWRDBUS_OUT[37]);
buf B_PPCMPLBWRDBUS38 (PPCMPLBWRDBUS[38], PPCMPLBWRDBUS_OUT[38]);
buf B_PPCMPLBWRDBUS39 (PPCMPLBWRDBUS[39], PPCMPLBWRDBUS_OUT[39]);
buf B_PPCMPLBWRDBUS40 (PPCMPLBWRDBUS[40], PPCMPLBWRDBUS_OUT[40]);
buf B_PPCMPLBWRDBUS41 (PPCMPLBWRDBUS[41], PPCMPLBWRDBUS_OUT[41]);
buf B_PPCMPLBWRDBUS42 (PPCMPLBWRDBUS[42], PPCMPLBWRDBUS_OUT[42]);
buf B_PPCMPLBWRDBUS43 (PPCMPLBWRDBUS[43], PPCMPLBWRDBUS_OUT[43]);
buf B_PPCMPLBWRDBUS44 (PPCMPLBWRDBUS[44], PPCMPLBWRDBUS_OUT[44]);
buf B_PPCMPLBWRDBUS45 (PPCMPLBWRDBUS[45], PPCMPLBWRDBUS_OUT[45]);
buf B_PPCMPLBWRDBUS46 (PPCMPLBWRDBUS[46], PPCMPLBWRDBUS_OUT[46]);
buf B_PPCMPLBWRDBUS47 (PPCMPLBWRDBUS[47], PPCMPLBWRDBUS_OUT[47]);
buf B_PPCMPLBWRDBUS48 (PPCMPLBWRDBUS[48], PPCMPLBWRDBUS_OUT[48]);
buf B_PPCMPLBWRDBUS49 (PPCMPLBWRDBUS[49], PPCMPLBWRDBUS_OUT[49]);
buf B_PPCMPLBWRDBUS50 (PPCMPLBWRDBUS[50], PPCMPLBWRDBUS_OUT[50]);
buf B_PPCMPLBWRDBUS51 (PPCMPLBWRDBUS[51], PPCMPLBWRDBUS_OUT[51]);
buf B_PPCMPLBWRDBUS52 (PPCMPLBWRDBUS[52], PPCMPLBWRDBUS_OUT[52]);
buf B_PPCMPLBWRDBUS53 (PPCMPLBWRDBUS[53], PPCMPLBWRDBUS_OUT[53]);
buf B_PPCMPLBWRDBUS54 (PPCMPLBWRDBUS[54], PPCMPLBWRDBUS_OUT[54]);
buf B_PPCMPLBWRDBUS55 (PPCMPLBWRDBUS[55], PPCMPLBWRDBUS_OUT[55]);
buf B_PPCMPLBWRDBUS56 (PPCMPLBWRDBUS[56], PPCMPLBWRDBUS_OUT[56]);
buf B_PPCMPLBWRDBUS57 (PPCMPLBWRDBUS[57], PPCMPLBWRDBUS_OUT[57]);
buf B_PPCMPLBWRDBUS58 (PPCMPLBWRDBUS[58], PPCMPLBWRDBUS_OUT[58]);
buf B_PPCMPLBWRDBUS59 (PPCMPLBWRDBUS[59], PPCMPLBWRDBUS_OUT[59]);
buf B_PPCMPLBWRDBUS60 (PPCMPLBWRDBUS[60], PPCMPLBWRDBUS_OUT[60]);
buf B_PPCMPLBWRDBUS61 (PPCMPLBWRDBUS[61], PPCMPLBWRDBUS_OUT[61]);
buf B_PPCMPLBWRDBUS62 (PPCMPLBWRDBUS[62], PPCMPLBWRDBUS_OUT[62]);
buf B_PPCMPLBWRDBUS63 (PPCMPLBWRDBUS[63], PPCMPLBWRDBUS_OUT[63]);
buf B_PPCMPLBWRDBUS64 (PPCMPLBWRDBUS[64], PPCMPLBWRDBUS_OUT[64]);
buf B_PPCMPLBWRDBUS65 (PPCMPLBWRDBUS[65], PPCMPLBWRDBUS_OUT[65]);
buf B_PPCMPLBWRDBUS66 (PPCMPLBWRDBUS[66], PPCMPLBWRDBUS_OUT[66]);
buf B_PPCMPLBWRDBUS67 (PPCMPLBWRDBUS[67], PPCMPLBWRDBUS_OUT[67]);
buf B_PPCMPLBWRDBUS68 (PPCMPLBWRDBUS[68], PPCMPLBWRDBUS_OUT[68]);
buf B_PPCMPLBWRDBUS69 (PPCMPLBWRDBUS[69], PPCMPLBWRDBUS_OUT[69]);
buf B_PPCMPLBWRDBUS70 (PPCMPLBWRDBUS[70], PPCMPLBWRDBUS_OUT[70]);
buf B_PPCMPLBWRDBUS71 (PPCMPLBWRDBUS[71], PPCMPLBWRDBUS_OUT[71]);
buf B_PPCMPLBWRDBUS72 (PPCMPLBWRDBUS[72], PPCMPLBWRDBUS_OUT[72]);
buf B_PPCMPLBWRDBUS73 (PPCMPLBWRDBUS[73], PPCMPLBWRDBUS_OUT[73]);
buf B_PPCMPLBWRDBUS74 (PPCMPLBWRDBUS[74], PPCMPLBWRDBUS_OUT[74]);
buf B_PPCMPLBWRDBUS75 (PPCMPLBWRDBUS[75], PPCMPLBWRDBUS_OUT[75]);
buf B_PPCMPLBWRDBUS76 (PPCMPLBWRDBUS[76], PPCMPLBWRDBUS_OUT[76]);
buf B_PPCMPLBWRDBUS77 (PPCMPLBWRDBUS[77], PPCMPLBWRDBUS_OUT[77]);
buf B_PPCMPLBWRDBUS78 (PPCMPLBWRDBUS[78], PPCMPLBWRDBUS_OUT[78]);
buf B_PPCMPLBWRDBUS79 (PPCMPLBWRDBUS[79], PPCMPLBWRDBUS_OUT[79]);
buf B_PPCMPLBWRDBUS80 (PPCMPLBWRDBUS[80], PPCMPLBWRDBUS_OUT[80]);
buf B_PPCMPLBWRDBUS81 (PPCMPLBWRDBUS[81], PPCMPLBWRDBUS_OUT[81]);
buf B_PPCMPLBWRDBUS82 (PPCMPLBWRDBUS[82], PPCMPLBWRDBUS_OUT[82]);
buf B_PPCMPLBWRDBUS83 (PPCMPLBWRDBUS[83], PPCMPLBWRDBUS_OUT[83]);
buf B_PPCMPLBWRDBUS84 (PPCMPLBWRDBUS[84], PPCMPLBWRDBUS_OUT[84]);
buf B_PPCMPLBWRDBUS85 (PPCMPLBWRDBUS[85], PPCMPLBWRDBUS_OUT[85]);
buf B_PPCMPLBWRDBUS86 (PPCMPLBWRDBUS[86], PPCMPLBWRDBUS_OUT[86]);
buf B_PPCMPLBWRDBUS87 (PPCMPLBWRDBUS[87], PPCMPLBWRDBUS_OUT[87]);
buf B_PPCMPLBWRDBUS88 (PPCMPLBWRDBUS[88], PPCMPLBWRDBUS_OUT[88]);
buf B_PPCMPLBWRDBUS89 (PPCMPLBWRDBUS[89], PPCMPLBWRDBUS_OUT[89]);
buf B_PPCMPLBWRDBUS90 (PPCMPLBWRDBUS[90], PPCMPLBWRDBUS_OUT[90]);
buf B_PPCMPLBWRDBUS91 (PPCMPLBWRDBUS[91], PPCMPLBWRDBUS_OUT[91]);
buf B_PPCMPLBWRDBUS92 (PPCMPLBWRDBUS[92], PPCMPLBWRDBUS_OUT[92]);
buf B_PPCMPLBWRDBUS93 (PPCMPLBWRDBUS[93], PPCMPLBWRDBUS_OUT[93]);
buf B_PPCMPLBWRDBUS94 (PPCMPLBWRDBUS[94], PPCMPLBWRDBUS_OUT[94]);
buf B_PPCMPLBWRDBUS95 (PPCMPLBWRDBUS[95], PPCMPLBWRDBUS_OUT[95]);
buf B_PPCMPLBWRDBUS96 (PPCMPLBWRDBUS[96], PPCMPLBWRDBUS_OUT[96]);
buf B_PPCMPLBWRDBUS97 (PPCMPLBWRDBUS[97], PPCMPLBWRDBUS_OUT[97]);
buf B_PPCMPLBWRDBUS98 (PPCMPLBWRDBUS[98], PPCMPLBWRDBUS_OUT[98]);
buf B_PPCMPLBWRDBUS99 (PPCMPLBWRDBUS[99], PPCMPLBWRDBUS_OUT[99]);
buf B_PPCMPLBWRDBUS100 (PPCMPLBWRDBUS[100], PPCMPLBWRDBUS_OUT[100]);
buf B_PPCMPLBWRDBUS101 (PPCMPLBWRDBUS[101], PPCMPLBWRDBUS_OUT[101]);
buf B_PPCMPLBWRDBUS102 (PPCMPLBWRDBUS[102], PPCMPLBWRDBUS_OUT[102]);
buf B_PPCMPLBWRDBUS103 (PPCMPLBWRDBUS[103], PPCMPLBWRDBUS_OUT[103]);
buf B_PPCMPLBWRDBUS104 (PPCMPLBWRDBUS[104], PPCMPLBWRDBUS_OUT[104]);
buf B_PPCMPLBWRDBUS105 (PPCMPLBWRDBUS[105], PPCMPLBWRDBUS_OUT[105]);
buf B_PPCMPLBWRDBUS106 (PPCMPLBWRDBUS[106], PPCMPLBWRDBUS_OUT[106]);
buf B_PPCMPLBWRDBUS107 (PPCMPLBWRDBUS[107], PPCMPLBWRDBUS_OUT[107]);
buf B_PPCMPLBWRDBUS108 (PPCMPLBWRDBUS[108], PPCMPLBWRDBUS_OUT[108]);
buf B_PPCMPLBWRDBUS109 (PPCMPLBWRDBUS[109], PPCMPLBWRDBUS_OUT[109]);
buf B_PPCMPLBWRDBUS110 (PPCMPLBWRDBUS[110], PPCMPLBWRDBUS_OUT[110]);
buf B_PPCMPLBWRDBUS111 (PPCMPLBWRDBUS[111], PPCMPLBWRDBUS_OUT[111]);
buf B_PPCMPLBWRDBUS112 (PPCMPLBWRDBUS[112], PPCMPLBWRDBUS_OUT[112]);
buf B_PPCMPLBWRDBUS113 (PPCMPLBWRDBUS[113], PPCMPLBWRDBUS_OUT[113]);
buf B_PPCMPLBWRDBUS114 (PPCMPLBWRDBUS[114], PPCMPLBWRDBUS_OUT[114]);
buf B_PPCMPLBWRDBUS115 (PPCMPLBWRDBUS[115], PPCMPLBWRDBUS_OUT[115]);
buf B_PPCMPLBWRDBUS116 (PPCMPLBWRDBUS[116], PPCMPLBWRDBUS_OUT[116]);
buf B_PPCMPLBWRDBUS117 (PPCMPLBWRDBUS[117], PPCMPLBWRDBUS_OUT[117]);
buf B_PPCMPLBWRDBUS118 (PPCMPLBWRDBUS[118], PPCMPLBWRDBUS_OUT[118]);
buf B_PPCMPLBWRDBUS119 (PPCMPLBWRDBUS[119], PPCMPLBWRDBUS_OUT[119]);
buf B_PPCMPLBWRDBUS120 (PPCMPLBWRDBUS[120], PPCMPLBWRDBUS_OUT[120]);
buf B_PPCMPLBWRDBUS121 (PPCMPLBWRDBUS[121], PPCMPLBWRDBUS_OUT[121]);
buf B_PPCMPLBWRDBUS122 (PPCMPLBWRDBUS[122], PPCMPLBWRDBUS_OUT[122]);
buf B_PPCMPLBWRDBUS123 (PPCMPLBWRDBUS[123], PPCMPLBWRDBUS_OUT[123]);
buf B_PPCMPLBWRDBUS124 (PPCMPLBWRDBUS[124], PPCMPLBWRDBUS_OUT[124]);
buf B_PPCMPLBWRDBUS125 (PPCMPLBWRDBUS[125], PPCMPLBWRDBUS_OUT[125]);
buf B_PPCMPLBWRDBUS126 (PPCMPLBWRDBUS[126], PPCMPLBWRDBUS_OUT[126]);
buf B_PPCMPLBWRDBUS127 (PPCMPLBWRDBUS[127], PPCMPLBWRDBUS_OUT[127]);
buf B_PPCS0PLBADDRACK (PPCS0PLBADDRACK, PPCS0PLBADDRACK_OUT);
buf B_PPCS0PLBMBUSY0 (PPCS0PLBMBUSY[0], PPCS0PLBMBUSY_OUT[0]);
buf B_PPCS0PLBMBUSY1 (PPCS0PLBMBUSY[1], PPCS0PLBMBUSY_OUT[1]);
buf B_PPCS0PLBMBUSY2 (PPCS0PLBMBUSY[2], PPCS0PLBMBUSY_OUT[2]);
buf B_PPCS0PLBMBUSY3 (PPCS0PLBMBUSY[3], PPCS0PLBMBUSY_OUT[3]);
buf B_PPCS0PLBMIRQ0 (PPCS0PLBMIRQ[0], PPCS0PLBMIRQ_OUT[0]);
buf B_PPCS0PLBMIRQ1 (PPCS0PLBMIRQ[1], PPCS0PLBMIRQ_OUT[1]);
buf B_PPCS0PLBMIRQ2 (PPCS0PLBMIRQ[2], PPCS0PLBMIRQ_OUT[2]);
buf B_PPCS0PLBMIRQ3 (PPCS0PLBMIRQ[3], PPCS0PLBMIRQ_OUT[3]);
buf B_PPCS0PLBMRDERR0 (PPCS0PLBMRDERR[0], PPCS0PLBMRDERR_OUT[0]);
buf B_PPCS0PLBMRDERR1 (PPCS0PLBMRDERR[1], PPCS0PLBMRDERR_OUT[1]);
buf B_PPCS0PLBMRDERR2 (PPCS0PLBMRDERR[2], PPCS0PLBMRDERR_OUT[2]);
buf B_PPCS0PLBMRDERR3 (PPCS0PLBMRDERR[3], PPCS0PLBMRDERR_OUT[3]);
buf B_PPCS0PLBMWRERR0 (PPCS0PLBMWRERR[0], PPCS0PLBMWRERR_OUT[0]);
buf B_PPCS0PLBMWRERR1 (PPCS0PLBMWRERR[1], PPCS0PLBMWRERR_OUT[1]);
buf B_PPCS0PLBMWRERR2 (PPCS0PLBMWRERR[2], PPCS0PLBMWRERR_OUT[2]);
buf B_PPCS0PLBMWRERR3 (PPCS0PLBMWRERR[3], PPCS0PLBMWRERR_OUT[3]);
buf B_PPCS0PLBRDBTERM (PPCS0PLBRDBTERM, PPCS0PLBRDBTERM_OUT);
buf B_PPCS0PLBRDCOMP (PPCS0PLBRDCOMP, PPCS0PLBRDCOMP_OUT);
buf B_PPCS0PLBRDDACK (PPCS0PLBRDDACK, PPCS0PLBRDDACK_OUT);
buf B_PPCS0PLBRDDBUS0 (PPCS0PLBRDDBUS[0], PPCS0PLBRDDBUS_OUT[0]);
buf B_PPCS0PLBRDDBUS1 (PPCS0PLBRDDBUS[1], PPCS0PLBRDDBUS_OUT[1]);
buf B_PPCS0PLBRDDBUS2 (PPCS0PLBRDDBUS[2], PPCS0PLBRDDBUS_OUT[2]);
buf B_PPCS0PLBRDDBUS3 (PPCS0PLBRDDBUS[3], PPCS0PLBRDDBUS_OUT[3]);
buf B_PPCS0PLBRDDBUS4 (PPCS0PLBRDDBUS[4], PPCS0PLBRDDBUS_OUT[4]);
buf B_PPCS0PLBRDDBUS5 (PPCS0PLBRDDBUS[5], PPCS0PLBRDDBUS_OUT[5]);
buf B_PPCS0PLBRDDBUS6 (PPCS0PLBRDDBUS[6], PPCS0PLBRDDBUS_OUT[6]);
buf B_PPCS0PLBRDDBUS7 (PPCS0PLBRDDBUS[7], PPCS0PLBRDDBUS_OUT[7]);
buf B_PPCS0PLBRDDBUS8 (PPCS0PLBRDDBUS[8], PPCS0PLBRDDBUS_OUT[8]);
buf B_PPCS0PLBRDDBUS9 (PPCS0PLBRDDBUS[9], PPCS0PLBRDDBUS_OUT[9]);
buf B_PPCS0PLBRDDBUS10 (PPCS0PLBRDDBUS[10], PPCS0PLBRDDBUS_OUT[10]);
buf B_PPCS0PLBRDDBUS11 (PPCS0PLBRDDBUS[11], PPCS0PLBRDDBUS_OUT[11]);
buf B_PPCS0PLBRDDBUS12 (PPCS0PLBRDDBUS[12], PPCS0PLBRDDBUS_OUT[12]);
buf B_PPCS0PLBRDDBUS13 (PPCS0PLBRDDBUS[13], PPCS0PLBRDDBUS_OUT[13]);
buf B_PPCS0PLBRDDBUS14 (PPCS0PLBRDDBUS[14], PPCS0PLBRDDBUS_OUT[14]);
buf B_PPCS0PLBRDDBUS15 (PPCS0PLBRDDBUS[15], PPCS0PLBRDDBUS_OUT[15]);
buf B_PPCS0PLBRDDBUS16 (PPCS0PLBRDDBUS[16], PPCS0PLBRDDBUS_OUT[16]);
buf B_PPCS0PLBRDDBUS17 (PPCS0PLBRDDBUS[17], PPCS0PLBRDDBUS_OUT[17]);
buf B_PPCS0PLBRDDBUS18 (PPCS0PLBRDDBUS[18], PPCS0PLBRDDBUS_OUT[18]);
buf B_PPCS0PLBRDDBUS19 (PPCS0PLBRDDBUS[19], PPCS0PLBRDDBUS_OUT[19]);
buf B_PPCS0PLBRDDBUS20 (PPCS0PLBRDDBUS[20], PPCS0PLBRDDBUS_OUT[20]);
buf B_PPCS0PLBRDDBUS21 (PPCS0PLBRDDBUS[21], PPCS0PLBRDDBUS_OUT[21]);
buf B_PPCS0PLBRDDBUS22 (PPCS0PLBRDDBUS[22], PPCS0PLBRDDBUS_OUT[22]);
buf B_PPCS0PLBRDDBUS23 (PPCS0PLBRDDBUS[23], PPCS0PLBRDDBUS_OUT[23]);
buf B_PPCS0PLBRDDBUS24 (PPCS0PLBRDDBUS[24], PPCS0PLBRDDBUS_OUT[24]);
buf B_PPCS0PLBRDDBUS25 (PPCS0PLBRDDBUS[25], PPCS0PLBRDDBUS_OUT[25]);
buf B_PPCS0PLBRDDBUS26 (PPCS0PLBRDDBUS[26], PPCS0PLBRDDBUS_OUT[26]);
buf B_PPCS0PLBRDDBUS27 (PPCS0PLBRDDBUS[27], PPCS0PLBRDDBUS_OUT[27]);
buf B_PPCS0PLBRDDBUS28 (PPCS0PLBRDDBUS[28], PPCS0PLBRDDBUS_OUT[28]);
buf B_PPCS0PLBRDDBUS29 (PPCS0PLBRDDBUS[29], PPCS0PLBRDDBUS_OUT[29]);
buf B_PPCS0PLBRDDBUS30 (PPCS0PLBRDDBUS[30], PPCS0PLBRDDBUS_OUT[30]);
buf B_PPCS0PLBRDDBUS31 (PPCS0PLBRDDBUS[31], PPCS0PLBRDDBUS_OUT[31]);
buf B_PPCS0PLBRDDBUS32 (PPCS0PLBRDDBUS[32], PPCS0PLBRDDBUS_OUT[32]);
buf B_PPCS0PLBRDDBUS33 (PPCS0PLBRDDBUS[33], PPCS0PLBRDDBUS_OUT[33]);
buf B_PPCS0PLBRDDBUS34 (PPCS0PLBRDDBUS[34], PPCS0PLBRDDBUS_OUT[34]);
buf B_PPCS0PLBRDDBUS35 (PPCS0PLBRDDBUS[35], PPCS0PLBRDDBUS_OUT[35]);
buf B_PPCS0PLBRDDBUS36 (PPCS0PLBRDDBUS[36], PPCS0PLBRDDBUS_OUT[36]);
buf B_PPCS0PLBRDDBUS37 (PPCS0PLBRDDBUS[37], PPCS0PLBRDDBUS_OUT[37]);
buf B_PPCS0PLBRDDBUS38 (PPCS0PLBRDDBUS[38], PPCS0PLBRDDBUS_OUT[38]);
buf B_PPCS0PLBRDDBUS39 (PPCS0PLBRDDBUS[39], PPCS0PLBRDDBUS_OUT[39]);
buf B_PPCS0PLBRDDBUS40 (PPCS0PLBRDDBUS[40], PPCS0PLBRDDBUS_OUT[40]);
buf B_PPCS0PLBRDDBUS41 (PPCS0PLBRDDBUS[41], PPCS0PLBRDDBUS_OUT[41]);
buf B_PPCS0PLBRDDBUS42 (PPCS0PLBRDDBUS[42], PPCS0PLBRDDBUS_OUT[42]);
buf B_PPCS0PLBRDDBUS43 (PPCS0PLBRDDBUS[43], PPCS0PLBRDDBUS_OUT[43]);
buf B_PPCS0PLBRDDBUS44 (PPCS0PLBRDDBUS[44], PPCS0PLBRDDBUS_OUT[44]);
buf B_PPCS0PLBRDDBUS45 (PPCS0PLBRDDBUS[45], PPCS0PLBRDDBUS_OUT[45]);
buf B_PPCS0PLBRDDBUS46 (PPCS0PLBRDDBUS[46], PPCS0PLBRDDBUS_OUT[46]);
buf B_PPCS0PLBRDDBUS47 (PPCS0PLBRDDBUS[47], PPCS0PLBRDDBUS_OUT[47]);
buf B_PPCS0PLBRDDBUS48 (PPCS0PLBRDDBUS[48], PPCS0PLBRDDBUS_OUT[48]);
buf B_PPCS0PLBRDDBUS49 (PPCS0PLBRDDBUS[49], PPCS0PLBRDDBUS_OUT[49]);
buf B_PPCS0PLBRDDBUS50 (PPCS0PLBRDDBUS[50], PPCS0PLBRDDBUS_OUT[50]);
buf B_PPCS0PLBRDDBUS51 (PPCS0PLBRDDBUS[51], PPCS0PLBRDDBUS_OUT[51]);
buf B_PPCS0PLBRDDBUS52 (PPCS0PLBRDDBUS[52], PPCS0PLBRDDBUS_OUT[52]);
buf B_PPCS0PLBRDDBUS53 (PPCS0PLBRDDBUS[53], PPCS0PLBRDDBUS_OUT[53]);
buf B_PPCS0PLBRDDBUS54 (PPCS0PLBRDDBUS[54], PPCS0PLBRDDBUS_OUT[54]);
buf B_PPCS0PLBRDDBUS55 (PPCS0PLBRDDBUS[55], PPCS0PLBRDDBUS_OUT[55]);
buf B_PPCS0PLBRDDBUS56 (PPCS0PLBRDDBUS[56], PPCS0PLBRDDBUS_OUT[56]);
buf B_PPCS0PLBRDDBUS57 (PPCS0PLBRDDBUS[57], PPCS0PLBRDDBUS_OUT[57]);
buf B_PPCS0PLBRDDBUS58 (PPCS0PLBRDDBUS[58], PPCS0PLBRDDBUS_OUT[58]);
buf B_PPCS0PLBRDDBUS59 (PPCS0PLBRDDBUS[59], PPCS0PLBRDDBUS_OUT[59]);
buf B_PPCS0PLBRDDBUS60 (PPCS0PLBRDDBUS[60], PPCS0PLBRDDBUS_OUT[60]);
buf B_PPCS0PLBRDDBUS61 (PPCS0PLBRDDBUS[61], PPCS0PLBRDDBUS_OUT[61]);
buf B_PPCS0PLBRDDBUS62 (PPCS0PLBRDDBUS[62], PPCS0PLBRDDBUS_OUT[62]);
buf B_PPCS0PLBRDDBUS63 (PPCS0PLBRDDBUS[63], PPCS0PLBRDDBUS_OUT[63]);
buf B_PPCS0PLBRDDBUS64 (PPCS0PLBRDDBUS[64], PPCS0PLBRDDBUS_OUT[64]);
buf B_PPCS0PLBRDDBUS65 (PPCS0PLBRDDBUS[65], PPCS0PLBRDDBUS_OUT[65]);
buf B_PPCS0PLBRDDBUS66 (PPCS0PLBRDDBUS[66], PPCS0PLBRDDBUS_OUT[66]);
buf B_PPCS0PLBRDDBUS67 (PPCS0PLBRDDBUS[67], PPCS0PLBRDDBUS_OUT[67]);
buf B_PPCS0PLBRDDBUS68 (PPCS0PLBRDDBUS[68], PPCS0PLBRDDBUS_OUT[68]);
buf B_PPCS0PLBRDDBUS69 (PPCS0PLBRDDBUS[69], PPCS0PLBRDDBUS_OUT[69]);
buf B_PPCS0PLBRDDBUS70 (PPCS0PLBRDDBUS[70], PPCS0PLBRDDBUS_OUT[70]);
buf B_PPCS0PLBRDDBUS71 (PPCS0PLBRDDBUS[71], PPCS0PLBRDDBUS_OUT[71]);
buf B_PPCS0PLBRDDBUS72 (PPCS0PLBRDDBUS[72], PPCS0PLBRDDBUS_OUT[72]);
buf B_PPCS0PLBRDDBUS73 (PPCS0PLBRDDBUS[73], PPCS0PLBRDDBUS_OUT[73]);
buf B_PPCS0PLBRDDBUS74 (PPCS0PLBRDDBUS[74], PPCS0PLBRDDBUS_OUT[74]);
buf B_PPCS0PLBRDDBUS75 (PPCS0PLBRDDBUS[75], PPCS0PLBRDDBUS_OUT[75]);
buf B_PPCS0PLBRDDBUS76 (PPCS0PLBRDDBUS[76], PPCS0PLBRDDBUS_OUT[76]);
buf B_PPCS0PLBRDDBUS77 (PPCS0PLBRDDBUS[77], PPCS0PLBRDDBUS_OUT[77]);
buf B_PPCS0PLBRDDBUS78 (PPCS0PLBRDDBUS[78], PPCS0PLBRDDBUS_OUT[78]);
buf B_PPCS0PLBRDDBUS79 (PPCS0PLBRDDBUS[79], PPCS0PLBRDDBUS_OUT[79]);
buf B_PPCS0PLBRDDBUS80 (PPCS0PLBRDDBUS[80], PPCS0PLBRDDBUS_OUT[80]);
buf B_PPCS0PLBRDDBUS81 (PPCS0PLBRDDBUS[81], PPCS0PLBRDDBUS_OUT[81]);
buf B_PPCS0PLBRDDBUS82 (PPCS0PLBRDDBUS[82], PPCS0PLBRDDBUS_OUT[82]);
buf B_PPCS0PLBRDDBUS83 (PPCS0PLBRDDBUS[83], PPCS0PLBRDDBUS_OUT[83]);
buf B_PPCS0PLBRDDBUS84 (PPCS0PLBRDDBUS[84], PPCS0PLBRDDBUS_OUT[84]);
buf B_PPCS0PLBRDDBUS85 (PPCS0PLBRDDBUS[85], PPCS0PLBRDDBUS_OUT[85]);
buf B_PPCS0PLBRDDBUS86 (PPCS0PLBRDDBUS[86], PPCS0PLBRDDBUS_OUT[86]);
buf B_PPCS0PLBRDDBUS87 (PPCS0PLBRDDBUS[87], PPCS0PLBRDDBUS_OUT[87]);
buf B_PPCS0PLBRDDBUS88 (PPCS0PLBRDDBUS[88], PPCS0PLBRDDBUS_OUT[88]);
buf B_PPCS0PLBRDDBUS89 (PPCS0PLBRDDBUS[89], PPCS0PLBRDDBUS_OUT[89]);
buf B_PPCS0PLBRDDBUS90 (PPCS0PLBRDDBUS[90], PPCS0PLBRDDBUS_OUT[90]);
buf B_PPCS0PLBRDDBUS91 (PPCS0PLBRDDBUS[91], PPCS0PLBRDDBUS_OUT[91]);
buf B_PPCS0PLBRDDBUS92 (PPCS0PLBRDDBUS[92], PPCS0PLBRDDBUS_OUT[92]);
buf B_PPCS0PLBRDDBUS93 (PPCS0PLBRDDBUS[93], PPCS0PLBRDDBUS_OUT[93]);
buf B_PPCS0PLBRDDBUS94 (PPCS0PLBRDDBUS[94], PPCS0PLBRDDBUS_OUT[94]);
buf B_PPCS0PLBRDDBUS95 (PPCS0PLBRDDBUS[95], PPCS0PLBRDDBUS_OUT[95]);
buf B_PPCS0PLBRDDBUS96 (PPCS0PLBRDDBUS[96], PPCS0PLBRDDBUS_OUT[96]);
buf B_PPCS0PLBRDDBUS97 (PPCS0PLBRDDBUS[97], PPCS0PLBRDDBUS_OUT[97]);
buf B_PPCS0PLBRDDBUS98 (PPCS0PLBRDDBUS[98], PPCS0PLBRDDBUS_OUT[98]);
buf B_PPCS0PLBRDDBUS99 (PPCS0PLBRDDBUS[99], PPCS0PLBRDDBUS_OUT[99]);
buf B_PPCS0PLBRDDBUS100 (PPCS0PLBRDDBUS[100], PPCS0PLBRDDBUS_OUT[100]);
buf B_PPCS0PLBRDDBUS101 (PPCS0PLBRDDBUS[101], PPCS0PLBRDDBUS_OUT[101]);
buf B_PPCS0PLBRDDBUS102 (PPCS0PLBRDDBUS[102], PPCS0PLBRDDBUS_OUT[102]);
buf B_PPCS0PLBRDDBUS103 (PPCS0PLBRDDBUS[103], PPCS0PLBRDDBUS_OUT[103]);
buf B_PPCS0PLBRDDBUS104 (PPCS0PLBRDDBUS[104], PPCS0PLBRDDBUS_OUT[104]);
buf B_PPCS0PLBRDDBUS105 (PPCS0PLBRDDBUS[105], PPCS0PLBRDDBUS_OUT[105]);
buf B_PPCS0PLBRDDBUS106 (PPCS0PLBRDDBUS[106], PPCS0PLBRDDBUS_OUT[106]);
buf B_PPCS0PLBRDDBUS107 (PPCS0PLBRDDBUS[107], PPCS0PLBRDDBUS_OUT[107]);
buf B_PPCS0PLBRDDBUS108 (PPCS0PLBRDDBUS[108], PPCS0PLBRDDBUS_OUT[108]);
buf B_PPCS0PLBRDDBUS109 (PPCS0PLBRDDBUS[109], PPCS0PLBRDDBUS_OUT[109]);
buf B_PPCS0PLBRDDBUS110 (PPCS0PLBRDDBUS[110], PPCS0PLBRDDBUS_OUT[110]);
buf B_PPCS0PLBRDDBUS111 (PPCS0PLBRDDBUS[111], PPCS0PLBRDDBUS_OUT[111]);
buf B_PPCS0PLBRDDBUS112 (PPCS0PLBRDDBUS[112], PPCS0PLBRDDBUS_OUT[112]);
buf B_PPCS0PLBRDDBUS113 (PPCS0PLBRDDBUS[113], PPCS0PLBRDDBUS_OUT[113]);
buf B_PPCS0PLBRDDBUS114 (PPCS0PLBRDDBUS[114], PPCS0PLBRDDBUS_OUT[114]);
buf B_PPCS0PLBRDDBUS115 (PPCS0PLBRDDBUS[115], PPCS0PLBRDDBUS_OUT[115]);
buf B_PPCS0PLBRDDBUS116 (PPCS0PLBRDDBUS[116], PPCS0PLBRDDBUS_OUT[116]);
buf B_PPCS0PLBRDDBUS117 (PPCS0PLBRDDBUS[117], PPCS0PLBRDDBUS_OUT[117]);
buf B_PPCS0PLBRDDBUS118 (PPCS0PLBRDDBUS[118], PPCS0PLBRDDBUS_OUT[118]);
buf B_PPCS0PLBRDDBUS119 (PPCS0PLBRDDBUS[119], PPCS0PLBRDDBUS_OUT[119]);
buf B_PPCS0PLBRDDBUS120 (PPCS0PLBRDDBUS[120], PPCS0PLBRDDBUS_OUT[120]);
buf B_PPCS0PLBRDDBUS121 (PPCS0PLBRDDBUS[121], PPCS0PLBRDDBUS_OUT[121]);
buf B_PPCS0PLBRDDBUS122 (PPCS0PLBRDDBUS[122], PPCS0PLBRDDBUS_OUT[122]);
buf B_PPCS0PLBRDDBUS123 (PPCS0PLBRDDBUS[123], PPCS0PLBRDDBUS_OUT[123]);
buf B_PPCS0PLBRDDBUS124 (PPCS0PLBRDDBUS[124], PPCS0PLBRDDBUS_OUT[124]);
buf B_PPCS0PLBRDDBUS125 (PPCS0PLBRDDBUS[125], PPCS0PLBRDDBUS_OUT[125]);
buf B_PPCS0PLBRDDBUS126 (PPCS0PLBRDDBUS[126], PPCS0PLBRDDBUS_OUT[126]);
buf B_PPCS0PLBRDDBUS127 (PPCS0PLBRDDBUS[127], PPCS0PLBRDDBUS_OUT[127]);
buf B_PPCS0PLBRDWDADDR0 (PPCS0PLBRDWDADDR[0], PPCS0PLBRDWDADDR_OUT[0]);
buf B_PPCS0PLBRDWDADDR1 (PPCS0PLBRDWDADDR[1], PPCS0PLBRDWDADDR_OUT[1]);
buf B_PPCS0PLBRDWDADDR2 (PPCS0PLBRDWDADDR[2], PPCS0PLBRDWDADDR_OUT[2]);
buf B_PPCS0PLBRDWDADDR3 (PPCS0PLBRDWDADDR[3], PPCS0PLBRDWDADDR_OUT[3]);
buf B_PPCS0PLBREARBITRATE (PPCS0PLBREARBITRATE, PPCS0PLBREARBITRATE_OUT);
buf B_PPCS0PLBSSIZE0 (PPCS0PLBSSIZE[0], PPCS0PLBSSIZE_OUT[0]);
buf B_PPCS0PLBSSIZE1 (PPCS0PLBSSIZE[1], PPCS0PLBSSIZE_OUT[1]);
buf B_PPCS0PLBWAIT (PPCS0PLBWAIT, PPCS0PLBWAIT_OUT);
buf B_PPCS0PLBWRBTERM (PPCS0PLBWRBTERM, PPCS0PLBWRBTERM_OUT);
buf B_PPCS0PLBWRCOMP (PPCS0PLBWRCOMP, PPCS0PLBWRCOMP_OUT);
buf B_PPCS0PLBWRDACK (PPCS0PLBWRDACK, PPCS0PLBWRDACK_OUT);
buf B_PPCS1PLBADDRACK (PPCS1PLBADDRACK, PPCS1PLBADDRACK_OUT);
buf B_PPCS1PLBMBUSY0 (PPCS1PLBMBUSY[0], PPCS1PLBMBUSY_OUT[0]);
buf B_PPCS1PLBMBUSY1 (PPCS1PLBMBUSY[1], PPCS1PLBMBUSY_OUT[1]);
buf B_PPCS1PLBMBUSY2 (PPCS1PLBMBUSY[2], PPCS1PLBMBUSY_OUT[2]);
buf B_PPCS1PLBMBUSY3 (PPCS1PLBMBUSY[3], PPCS1PLBMBUSY_OUT[3]);
buf B_PPCS1PLBMIRQ0 (PPCS1PLBMIRQ[0], PPCS1PLBMIRQ_OUT[0]);
buf B_PPCS1PLBMIRQ1 (PPCS1PLBMIRQ[1], PPCS1PLBMIRQ_OUT[1]);
buf B_PPCS1PLBMIRQ2 (PPCS1PLBMIRQ[2], PPCS1PLBMIRQ_OUT[2]);
buf B_PPCS1PLBMIRQ3 (PPCS1PLBMIRQ[3], PPCS1PLBMIRQ_OUT[3]);
buf B_PPCS1PLBMRDERR0 (PPCS1PLBMRDERR[0], PPCS1PLBMRDERR_OUT[0]);
buf B_PPCS1PLBMRDERR1 (PPCS1PLBMRDERR[1], PPCS1PLBMRDERR_OUT[1]);
buf B_PPCS1PLBMRDERR2 (PPCS1PLBMRDERR[2], PPCS1PLBMRDERR_OUT[2]);
buf B_PPCS1PLBMRDERR3 (PPCS1PLBMRDERR[3], PPCS1PLBMRDERR_OUT[3]);
buf B_PPCS1PLBMWRERR0 (PPCS1PLBMWRERR[0], PPCS1PLBMWRERR_OUT[0]);
buf B_PPCS1PLBMWRERR1 (PPCS1PLBMWRERR[1], PPCS1PLBMWRERR_OUT[1]);
buf B_PPCS1PLBMWRERR2 (PPCS1PLBMWRERR[2], PPCS1PLBMWRERR_OUT[2]);
buf B_PPCS1PLBMWRERR3 (PPCS1PLBMWRERR[3], PPCS1PLBMWRERR_OUT[3]);
buf B_PPCS1PLBRDBTERM (PPCS1PLBRDBTERM, PPCS1PLBRDBTERM_OUT);
buf B_PPCS1PLBRDCOMP (PPCS1PLBRDCOMP, PPCS1PLBRDCOMP_OUT);
buf B_PPCS1PLBRDDACK (PPCS1PLBRDDACK, PPCS1PLBRDDACK_OUT);
buf B_PPCS1PLBRDDBUS0 (PPCS1PLBRDDBUS[0], PPCS1PLBRDDBUS_OUT[0]);
buf B_PPCS1PLBRDDBUS1 (PPCS1PLBRDDBUS[1], PPCS1PLBRDDBUS_OUT[1]);
buf B_PPCS1PLBRDDBUS2 (PPCS1PLBRDDBUS[2], PPCS1PLBRDDBUS_OUT[2]);
buf B_PPCS1PLBRDDBUS3 (PPCS1PLBRDDBUS[3], PPCS1PLBRDDBUS_OUT[3]);
buf B_PPCS1PLBRDDBUS4 (PPCS1PLBRDDBUS[4], PPCS1PLBRDDBUS_OUT[4]);
buf B_PPCS1PLBRDDBUS5 (PPCS1PLBRDDBUS[5], PPCS1PLBRDDBUS_OUT[5]);
buf B_PPCS1PLBRDDBUS6 (PPCS1PLBRDDBUS[6], PPCS1PLBRDDBUS_OUT[6]);
buf B_PPCS1PLBRDDBUS7 (PPCS1PLBRDDBUS[7], PPCS1PLBRDDBUS_OUT[7]);
buf B_PPCS1PLBRDDBUS8 (PPCS1PLBRDDBUS[8], PPCS1PLBRDDBUS_OUT[8]);
buf B_PPCS1PLBRDDBUS9 (PPCS1PLBRDDBUS[9], PPCS1PLBRDDBUS_OUT[9]);
buf B_PPCS1PLBRDDBUS10 (PPCS1PLBRDDBUS[10], PPCS1PLBRDDBUS_OUT[10]);
buf B_PPCS1PLBRDDBUS11 (PPCS1PLBRDDBUS[11], PPCS1PLBRDDBUS_OUT[11]);
buf B_PPCS1PLBRDDBUS12 (PPCS1PLBRDDBUS[12], PPCS1PLBRDDBUS_OUT[12]);
buf B_PPCS1PLBRDDBUS13 (PPCS1PLBRDDBUS[13], PPCS1PLBRDDBUS_OUT[13]);
buf B_PPCS1PLBRDDBUS14 (PPCS1PLBRDDBUS[14], PPCS1PLBRDDBUS_OUT[14]);
buf B_PPCS1PLBRDDBUS15 (PPCS1PLBRDDBUS[15], PPCS1PLBRDDBUS_OUT[15]);
buf B_PPCS1PLBRDDBUS16 (PPCS1PLBRDDBUS[16], PPCS1PLBRDDBUS_OUT[16]);
buf B_PPCS1PLBRDDBUS17 (PPCS1PLBRDDBUS[17], PPCS1PLBRDDBUS_OUT[17]);
buf B_PPCS1PLBRDDBUS18 (PPCS1PLBRDDBUS[18], PPCS1PLBRDDBUS_OUT[18]);
buf B_PPCS1PLBRDDBUS19 (PPCS1PLBRDDBUS[19], PPCS1PLBRDDBUS_OUT[19]);
buf B_PPCS1PLBRDDBUS20 (PPCS1PLBRDDBUS[20], PPCS1PLBRDDBUS_OUT[20]);
buf B_PPCS1PLBRDDBUS21 (PPCS1PLBRDDBUS[21], PPCS1PLBRDDBUS_OUT[21]);
buf B_PPCS1PLBRDDBUS22 (PPCS1PLBRDDBUS[22], PPCS1PLBRDDBUS_OUT[22]);
buf B_PPCS1PLBRDDBUS23 (PPCS1PLBRDDBUS[23], PPCS1PLBRDDBUS_OUT[23]);
buf B_PPCS1PLBRDDBUS24 (PPCS1PLBRDDBUS[24], PPCS1PLBRDDBUS_OUT[24]);
buf B_PPCS1PLBRDDBUS25 (PPCS1PLBRDDBUS[25], PPCS1PLBRDDBUS_OUT[25]);
buf B_PPCS1PLBRDDBUS26 (PPCS1PLBRDDBUS[26], PPCS1PLBRDDBUS_OUT[26]);
buf B_PPCS1PLBRDDBUS27 (PPCS1PLBRDDBUS[27], PPCS1PLBRDDBUS_OUT[27]);
buf B_PPCS1PLBRDDBUS28 (PPCS1PLBRDDBUS[28], PPCS1PLBRDDBUS_OUT[28]);
buf B_PPCS1PLBRDDBUS29 (PPCS1PLBRDDBUS[29], PPCS1PLBRDDBUS_OUT[29]);
buf B_PPCS1PLBRDDBUS30 (PPCS1PLBRDDBUS[30], PPCS1PLBRDDBUS_OUT[30]);
buf B_PPCS1PLBRDDBUS31 (PPCS1PLBRDDBUS[31], PPCS1PLBRDDBUS_OUT[31]);
buf B_PPCS1PLBRDDBUS32 (PPCS1PLBRDDBUS[32], PPCS1PLBRDDBUS_OUT[32]);
buf B_PPCS1PLBRDDBUS33 (PPCS1PLBRDDBUS[33], PPCS1PLBRDDBUS_OUT[33]);
buf B_PPCS1PLBRDDBUS34 (PPCS1PLBRDDBUS[34], PPCS1PLBRDDBUS_OUT[34]);
buf B_PPCS1PLBRDDBUS35 (PPCS1PLBRDDBUS[35], PPCS1PLBRDDBUS_OUT[35]);
buf B_PPCS1PLBRDDBUS36 (PPCS1PLBRDDBUS[36], PPCS1PLBRDDBUS_OUT[36]);
buf B_PPCS1PLBRDDBUS37 (PPCS1PLBRDDBUS[37], PPCS1PLBRDDBUS_OUT[37]);
buf B_PPCS1PLBRDDBUS38 (PPCS1PLBRDDBUS[38], PPCS1PLBRDDBUS_OUT[38]);
buf B_PPCS1PLBRDDBUS39 (PPCS1PLBRDDBUS[39], PPCS1PLBRDDBUS_OUT[39]);
buf B_PPCS1PLBRDDBUS40 (PPCS1PLBRDDBUS[40], PPCS1PLBRDDBUS_OUT[40]);
buf B_PPCS1PLBRDDBUS41 (PPCS1PLBRDDBUS[41], PPCS1PLBRDDBUS_OUT[41]);
buf B_PPCS1PLBRDDBUS42 (PPCS1PLBRDDBUS[42], PPCS1PLBRDDBUS_OUT[42]);
buf B_PPCS1PLBRDDBUS43 (PPCS1PLBRDDBUS[43], PPCS1PLBRDDBUS_OUT[43]);
buf B_PPCS1PLBRDDBUS44 (PPCS1PLBRDDBUS[44], PPCS1PLBRDDBUS_OUT[44]);
buf B_PPCS1PLBRDDBUS45 (PPCS1PLBRDDBUS[45], PPCS1PLBRDDBUS_OUT[45]);
buf B_PPCS1PLBRDDBUS46 (PPCS1PLBRDDBUS[46], PPCS1PLBRDDBUS_OUT[46]);
buf B_PPCS1PLBRDDBUS47 (PPCS1PLBRDDBUS[47], PPCS1PLBRDDBUS_OUT[47]);
buf B_PPCS1PLBRDDBUS48 (PPCS1PLBRDDBUS[48], PPCS1PLBRDDBUS_OUT[48]);
buf B_PPCS1PLBRDDBUS49 (PPCS1PLBRDDBUS[49], PPCS1PLBRDDBUS_OUT[49]);
buf B_PPCS1PLBRDDBUS50 (PPCS1PLBRDDBUS[50], PPCS1PLBRDDBUS_OUT[50]);
buf B_PPCS1PLBRDDBUS51 (PPCS1PLBRDDBUS[51], PPCS1PLBRDDBUS_OUT[51]);
buf B_PPCS1PLBRDDBUS52 (PPCS1PLBRDDBUS[52], PPCS1PLBRDDBUS_OUT[52]);
buf B_PPCS1PLBRDDBUS53 (PPCS1PLBRDDBUS[53], PPCS1PLBRDDBUS_OUT[53]);
buf B_PPCS1PLBRDDBUS54 (PPCS1PLBRDDBUS[54], PPCS1PLBRDDBUS_OUT[54]);
buf B_PPCS1PLBRDDBUS55 (PPCS1PLBRDDBUS[55], PPCS1PLBRDDBUS_OUT[55]);
buf B_PPCS1PLBRDDBUS56 (PPCS1PLBRDDBUS[56], PPCS1PLBRDDBUS_OUT[56]);
buf B_PPCS1PLBRDDBUS57 (PPCS1PLBRDDBUS[57], PPCS1PLBRDDBUS_OUT[57]);
buf B_PPCS1PLBRDDBUS58 (PPCS1PLBRDDBUS[58], PPCS1PLBRDDBUS_OUT[58]);
buf B_PPCS1PLBRDDBUS59 (PPCS1PLBRDDBUS[59], PPCS1PLBRDDBUS_OUT[59]);
buf B_PPCS1PLBRDDBUS60 (PPCS1PLBRDDBUS[60], PPCS1PLBRDDBUS_OUT[60]);
buf B_PPCS1PLBRDDBUS61 (PPCS1PLBRDDBUS[61], PPCS1PLBRDDBUS_OUT[61]);
buf B_PPCS1PLBRDDBUS62 (PPCS1PLBRDDBUS[62], PPCS1PLBRDDBUS_OUT[62]);
buf B_PPCS1PLBRDDBUS63 (PPCS1PLBRDDBUS[63], PPCS1PLBRDDBUS_OUT[63]);
buf B_PPCS1PLBRDDBUS64 (PPCS1PLBRDDBUS[64], PPCS1PLBRDDBUS_OUT[64]);
buf B_PPCS1PLBRDDBUS65 (PPCS1PLBRDDBUS[65], PPCS1PLBRDDBUS_OUT[65]);
buf B_PPCS1PLBRDDBUS66 (PPCS1PLBRDDBUS[66], PPCS1PLBRDDBUS_OUT[66]);
buf B_PPCS1PLBRDDBUS67 (PPCS1PLBRDDBUS[67], PPCS1PLBRDDBUS_OUT[67]);
buf B_PPCS1PLBRDDBUS68 (PPCS1PLBRDDBUS[68], PPCS1PLBRDDBUS_OUT[68]);
buf B_PPCS1PLBRDDBUS69 (PPCS1PLBRDDBUS[69], PPCS1PLBRDDBUS_OUT[69]);
buf B_PPCS1PLBRDDBUS70 (PPCS1PLBRDDBUS[70], PPCS1PLBRDDBUS_OUT[70]);
buf B_PPCS1PLBRDDBUS71 (PPCS1PLBRDDBUS[71], PPCS1PLBRDDBUS_OUT[71]);
buf B_PPCS1PLBRDDBUS72 (PPCS1PLBRDDBUS[72], PPCS1PLBRDDBUS_OUT[72]);
buf B_PPCS1PLBRDDBUS73 (PPCS1PLBRDDBUS[73], PPCS1PLBRDDBUS_OUT[73]);
buf B_PPCS1PLBRDDBUS74 (PPCS1PLBRDDBUS[74], PPCS1PLBRDDBUS_OUT[74]);
buf B_PPCS1PLBRDDBUS75 (PPCS1PLBRDDBUS[75], PPCS1PLBRDDBUS_OUT[75]);
buf B_PPCS1PLBRDDBUS76 (PPCS1PLBRDDBUS[76], PPCS1PLBRDDBUS_OUT[76]);
buf B_PPCS1PLBRDDBUS77 (PPCS1PLBRDDBUS[77], PPCS1PLBRDDBUS_OUT[77]);
buf B_PPCS1PLBRDDBUS78 (PPCS1PLBRDDBUS[78], PPCS1PLBRDDBUS_OUT[78]);
buf B_PPCS1PLBRDDBUS79 (PPCS1PLBRDDBUS[79], PPCS1PLBRDDBUS_OUT[79]);
buf B_PPCS1PLBRDDBUS80 (PPCS1PLBRDDBUS[80], PPCS1PLBRDDBUS_OUT[80]);
buf B_PPCS1PLBRDDBUS81 (PPCS1PLBRDDBUS[81], PPCS1PLBRDDBUS_OUT[81]);
buf B_PPCS1PLBRDDBUS82 (PPCS1PLBRDDBUS[82], PPCS1PLBRDDBUS_OUT[82]);
buf B_PPCS1PLBRDDBUS83 (PPCS1PLBRDDBUS[83], PPCS1PLBRDDBUS_OUT[83]);
buf B_PPCS1PLBRDDBUS84 (PPCS1PLBRDDBUS[84], PPCS1PLBRDDBUS_OUT[84]);
buf B_PPCS1PLBRDDBUS85 (PPCS1PLBRDDBUS[85], PPCS1PLBRDDBUS_OUT[85]);
buf B_PPCS1PLBRDDBUS86 (PPCS1PLBRDDBUS[86], PPCS1PLBRDDBUS_OUT[86]);
buf B_PPCS1PLBRDDBUS87 (PPCS1PLBRDDBUS[87], PPCS1PLBRDDBUS_OUT[87]);
buf B_PPCS1PLBRDDBUS88 (PPCS1PLBRDDBUS[88], PPCS1PLBRDDBUS_OUT[88]);
buf B_PPCS1PLBRDDBUS89 (PPCS1PLBRDDBUS[89], PPCS1PLBRDDBUS_OUT[89]);
buf B_PPCS1PLBRDDBUS90 (PPCS1PLBRDDBUS[90], PPCS1PLBRDDBUS_OUT[90]);
buf B_PPCS1PLBRDDBUS91 (PPCS1PLBRDDBUS[91], PPCS1PLBRDDBUS_OUT[91]);
buf B_PPCS1PLBRDDBUS92 (PPCS1PLBRDDBUS[92], PPCS1PLBRDDBUS_OUT[92]);
buf B_PPCS1PLBRDDBUS93 (PPCS1PLBRDDBUS[93], PPCS1PLBRDDBUS_OUT[93]);
buf B_PPCS1PLBRDDBUS94 (PPCS1PLBRDDBUS[94], PPCS1PLBRDDBUS_OUT[94]);
buf B_PPCS1PLBRDDBUS95 (PPCS1PLBRDDBUS[95], PPCS1PLBRDDBUS_OUT[95]);
buf B_PPCS1PLBRDDBUS96 (PPCS1PLBRDDBUS[96], PPCS1PLBRDDBUS_OUT[96]);
buf B_PPCS1PLBRDDBUS97 (PPCS1PLBRDDBUS[97], PPCS1PLBRDDBUS_OUT[97]);
buf B_PPCS1PLBRDDBUS98 (PPCS1PLBRDDBUS[98], PPCS1PLBRDDBUS_OUT[98]);
buf B_PPCS1PLBRDDBUS99 (PPCS1PLBRDDBUS[99], PPCS1PLBRDDBUS_OUT[99]);
buf B_PPCS1PLBRDDBUS100 (PPCS1PLBRDDBUS[100], PPCS1PLBRDDBUS_OUT[100]);
buf B_PPCS1PLBRDDBUS101 (PPCS1PLBRDDBUS[101], PPCS1PLBRDDBUS_OUT[101]);
buf B_PPCS1PLBRDDBUS102 (PPCS1PLBRDDBUS[102], PPCS1PLBRDDBUS_OUT[102]);
buf B_PPCS1PLBRDDBUS103 (PPCS1PLBRDDBUS[103], PPCS1PLBRDDBUS_OUT[103]);
buf B_PPCS1PLBRDDBUS104 (PPCS1PLBRDDBUS[104], PPCS1PLBRDDBUS_OUT[104]);
buf B_PPCS1PLBRDDBUS105 (PPCS1PLBRDDBUS[105], PPCS1PLBRDDBUS_OUT[105]);
buf B_PPCS1PLBRDDBUS106 (PPCS1PLBRDDBUS[106], PPCS1PLBRDDBUS_OUT[106]);
buf B_PPCS1PLBRDDBUS107 (PPCS1PLBRDDBUS[107], PPCS1PLBRDDBUS_OUT[107]);
buf B_PPCS1PLBRDDBUS108 (PPCS1PLBRDDBUS[108], PPCS1PLBRDDBUS_OUT[108]);
buf B_PPCS1PLBRDDBUS109 (PPCS1PLBRDDBUS[109], PPCS1PLBRDDBUS_OUT[109]);
buf B_PPCS1PLBRDDBUS110 (PPCS1PLBRDDBUS[110], PPCS1PLBRDDBUS_OUT[110]);
buf B_PPCS1PLBRDDBUS111 (PPCS1PLBRDDBUS[111], PPCS1PLBRDDBUS_OUT[111]);
buf B_PPCS1PLBRDDBUS112 (PPCS1PLBRDDBUS[112], PPCS1PLBRDDBUS_OUT[112]);
buf B_PPCS1PLBRDDBUS113 (PPCS1PLBRDDBUS[113], PPCS1PLBRDDBUS_OUT[113]);
buf B_PPCS1PLBRDDBUS114 (PPCS1PLBRDDBUS[114], PPCS1PLBRDDBUS_OUT[114]);
buf B_PPCS1PLBRDDBUS115 (PPCS1PLBRDDBUS[115], PPCS1PLBRDDBUS_OUT[115]);
buf B_PPCS1PLBRDDBUS116 (PPCS1PLBRDDBUS[116], PPCS1PLBRDDBUS_OUT[116]);
buf B_PPCS1PLBRDDBUS117 (PPCS1PLBRDDBUS[117], PPCS1PLBRDDBUS_OUT[117]);
buf B_PPCS1PLBRDDBUS118 (PPCS1PLBRDDBUS[118], PPCS1PLBRDDBUS_OUT[118]);
buf B_PPCS1PLBRDDBUS119 (PPCS1PLBRDDBUS[119], PPCS1PLBRDDBUS_OUT[119]);
buf B_PPCS1PLBRDDBUS120 (PPCS1PLBRDDBUS[120], PPCS1PLBRDDBUS_OUT[120]);
buf B_PPCS1PLBRDDBUS121 (PPCS1PLBRDDBUS[121], PPCS1PLBRDDBUS_OUT[121]);
buf B_PPCS1PLBRDDBUS122 (PPCS1PLBRDDBUS[122], PPCS1PLBRDDBUS_OUT[122]);
buf B_PPCS1PLBRDDBUS123 (PPCS1PLBRDDBUS[123], PPCS1PLBRDDBUS_OUT[123]);
buf B_PPCS1PLBRDDBUS124 (PPCS1PLBRDDBUS[124], PPCS1PLBRDDBUS_OUT[124]);
buf B_PPCS1PLBRDDBUS125 (PPCS1PLBRDDBUS[125], PPCS1PLBRDDBUS_OUT[125]);
buf B_PPCS1PLBRDDBUS126 (PPCS1PLBRDDBUS[126], PPCS1PLBRDDBUS_OUT[126]);
buf B_PPCS1PLBRDDBUS127 (PPCS1PLBRDDBUS[127], PPCS1PLBRDDBUS_OUT[127]);
buf B_PPCS1PLBRDWDADDR0 (PPCS1PLBRDWDADDR[0], PPCS1PLBRDWDADDR_OUT[0]);
buf B_PPCS1PLBRDWDADDR1 (PPCS1PLBRDWDADDR[1], PPCS1PLBRDWDADDR_OUT[1]);
buf B_PPCS1PLBRDWDADDR2 (PPCS1PLBRDWDADDR[2], PPCS1PLBRDWDADDR_OUT[2]);
buf B_PPCS1PLBRDWDADDR3 (PPCS1PLBRDWDADDR[3], PPCS1PLBRDWDADDR_OUT[3]);
buf B_PPCS1PLBREARBITRATE (PPCS1PLBREARBITRATE, PPCS1PLBREARBITRATE_OUT);
buf B_PPCS1PLBSSIZE0 (PPCS1PLBSSIZE[0], PPCS1PLBSSIZE_OUT[0]);
buf B_PPCS1PLBSSIZE1 (PPCS1PLBSSIZE[1], PPCS1PLBSSIZE_OUT[1]);
buf B_PPCS1PLBWAIT (PPCS1PLBWAIT, PPCS1PLBWAIT_OUT);
buf B_PPCS1PLBWRBTERM (PPCS1PLBWRBTERM, PPCS1PLBWRBTERM_OUT);
buf B_PPCS1PLBWRCOMP (PPCS1PLBWRCOMP, PPCS1PLBWRCOMP_OUT);
buf B_PPCS1PLBWRDACK (PPCS1PLBWRDACK, PPCS1PLBWRDACK_OUT);
buf B_APUFCMDECFPUOP (APUFCMDECFPUOP, APUFCMDECFPUOP_OUT);
buf B_APUFCMDECLDSTXFERSIZE0 (APUFCMDECLDSTXFERSIZE[0], APUFCMDECLDSTXFERSIZE_OUT[0]);
buf B_APUFCMDECLDSTXFERSIZE1 (APUFCMDECLDSTXFERSIZE[1], APUFCMDECLDSTXFERSIZE_OUT[1]);
buf B_APUFCMDECLDSTXFERSIZE2 (APUFCMDECLDSTXFERSIZE[2], APUFCMDECLDSTXFERSIZE_OUT[2]);
buf B_APUFCMDECLOAD (APUFCMDECLOAD, APUFCMDECLOAD_OUT);
buf B_APUFCMDECNONAUTON (APUFCMDECNONAUTON, APUFCMDECNONAUTON_OUT);
buf B_APUFCMDECSTORE (APUFCMDECSTORE, APUFCMDECSTORE_OUT);
buf B_APUFCMDECUDI0 (APUFCMDECUDI[0], APUFCMDECUDI_OUT[0]);
buf B_APUFCMDECUDI1 (APUFCMDECUDI[1], APUFCMDECUDI_OUT[1]);
buf B_APUFCMDECUDI2 (APUFCMDECUDI[2], APUFCMDECUDI_OUT[2]);
buf B_APUFCMDECUDI3 (APUFCMDECUDI[3], APUFCMDECUDI_OUT[3]);
buf B_APUFCMDECUDIVALID (APUFCMDECUDIVALID, APUFCMDECUDIVALID_OUT);
buf B_APUFCMENDIAN (APUFCMENDIAN, APUFCMENDIAN_OUT);
buf B_APUFCMFLUSH (APUFCMFLUSH, APUFCMFLUSH_OUT);
buf B_APUFCMINSTRUCTION0 (APUFCMINSTRUCTION[0], APUFCMINSTRUCTION_OUT[0]);
buf B_APUFCMINSTRUCTION1 (APUFCMINSTRUCTION[1], APUFCMINSTRUCTION_OUT[1]);
buf B_APUFCMINSTRUCTION2 (APUFCMINSTRUCTION[2], APUFCMINSTRUCTION_OUT[2]);
buf B_APUFCMINSTRUCTION3 (APUFCMINSTRUCTION[3], APUFCMINSTRUCTION_OUT[3]);
buf B_APUFCMINSTRUCTION4 (APUFCMINSTRUCTION[4], APUFCMINSTRUCTION_OUT[4]);
buf B_APUFCMINSTRUCTION5 (APUFCMINSTRUCTION[5], APUFCMINSTRUCTION_OUT[5]);
buf B_APUFCMINSTRUCTION6 (APUFCMINSTRUCTION[6], APUFCMINSTRUCTION_OUT[6]);
buf B_APUFCMINSTRUCTION7 (APUFCMINSTRUCTION[7], APUFCMINSTRUCTION_OUT[7]);
buf B_APUFCMINSTRUCTION8 (APUFCMINSTRUCTION[8], APUFCMINSTRUCTION_OUT[8]);
buf B_APUFCMINSTRUCTION9 (APUFCMINSTRUCTION[9], APUFCMINSTRUCTION_OUT[9]);
buf B_APUFCMINSTRUCTION10 (APUFCMINSTRUCTION[10], APUFCMINSTRUCTION_OUT[10]);
buf B_APUFCMINSTRUCTION11 (APUFCMINSTRUCTION[11], APUFCMINSTRUCTION_OUT[11]);
buf B_APUFCMINSTRUCTION12 (APUFCMINSTRUCTION[12], APUFCMINSTRUCTION_OUT[12]);
buf B_APUFCMINSTRUCTION13 (APUFCMINSTRUCTION[13], APUFCMINSTRUCTION_OUT[13]);
buf B_APUFCMINSTRUCTION14 (APUFCMINSTRUCTION[14], APUFCMINSTRUCTION_OUT[14]);
buf B_APUFCMINSTRUCTION15 (APUFCMINSTRUCTION[15], APUFCMINSTRUCTION_OUT[15]);
buf B_APUFCMINSTRUCTION16 (APUFCMINSTRUCTION[16], APUFCMINSTRUCTION_OUT[16]);
buf B_APUFCMINSTRUCTION17 (APUFCMINSTRUCTION[17], APUFCMINSTRUCTION_OUT[17]);
buf B_APUFCMINSTRUCTION18 (APUFCMINSTRUCTION[18], APUFCMINSTRUCTION_OUT[18]);
buf B_APUFCMINSTRUCTION19 (APUFCMINSTRUCTION[19], APUFCMINSTRUCTION_OUT[19]);
buf B_APUFCMINSTRUCTION20 (APUFCMINSTRUCTION[20], APUFCMINSTRUCTION_OUT[20]);
buf B_APUFCMINSTRUCTION21 (APUFCMINSTRUCTION[21], APUFCMINSTRUCTION_OUT[21]);
buf B_APUFCMINSTRUCTION22 (APUFCMINSTRUCTION[22], APUFCMINSTRUCTION_OUT[22]);
buf B_APUFCMINSTRUCTION23 (APUFCMINSTRUCTION[23], APUFCMINSTRUCTION_OUT[23]);
buf B_APUFCMINSTRUCTION24 (APUFCMINSTRUCTION[24], APUFCMINSTRUCTION_OUT[24]);
buf B_APUFCMINSTRUCTION25 (APUFCMINSTRUCTION[25], APUFCMINSTRUCTION_OUT[25]);
buf B_APUFCMINSTRUCTION26 (APUFCMINSTRUCTION[26], APUFCMINSTRUCTION_OUT[26]);
buf B_APUFCMINSTRUCTION27 (APUFCMINSTRUCTION[27], APUFCMINSTRUCTION_OUT[27]);
buf B_APUFCMINSTRUCTION28 (APUFCMINSTRUCTION[28], APUFCMINSTRUCTION_OUT[28]);
buf B_APUFCMINSTRUCTION29 (APUFCMINSTRUCTION[29], APUFCMINSTRUCTION_OUT[29]);
buf B_APUFCMINSTRUCTION30 (APUFCMINSTRUCTION[30], APUFCMINSTRUCTION_OUT[30]);
buf B_APUFCMINSTRUCTION31 (APUFCMINSTRUCTION[31], APUFCMINSTRUCTION_OUT[31]);
buf B_APUFCMINSTRVALID (APUFCMINSTRVALID, APUFCMINSTRVALID_OUT);
buf B_APUFCMLOADBYTEADDR0 (APUFCMLOADBYTEADDR[0], APUFCMLOADBYTEADDR_OUT[0]);
buf B_APUFCMLOADBYTEADDR1 (APUFCMLOADBYTEADDR[1], APUFCMLOADBYTEADDR_OUT[1]);
buf B_APUFCMLOADBYTEADDR2 (APUFCMLOADBYTEADDR[2], APUFCMLOADBYTEADDR_OUT[2]);
buf B_APUFCMLOADBYTEADDR3 (APUFCMLOADBYTEADDR[3], APUFCMLOADBYTEADDR_OUT[3]);
buf B_APUFCMLOADDATA0 (APUFCMLOADDATA[0], APUFCMLOADDATA_OUT[0]);
buf B_APUFCMLOADDATA1 (APUFCMLOADDATA[1], APUFCMLOADDATA_OUT[1]);
buf B_APUFCMLOADDATA2 (APUFCMLOADDATA[2], APUFCMLOADDATA_OUT[2]);
buf B_APUFCMLOADDATA3 (APUFCMLOADDATA[3], APUFCMLOADDATA_OUT[3]);
buf B_APUFCMLOADDATA4 (APUFCMLOADDATA[4], APUFCMLOADDATA_OUT[4]);
buf B_APUFCMLOADDATA5 (APUFCMLOADDATA[5], APUFCMLOADDATA_OUT[5]);
buf B_APUFCMLOADDATA6 (APUFCMLOADDATA[6], APUFCMLOADDATA_OUT[6]);
buf B_APUFCMLOADDATA7 (APUFCMLOADDATA[7], APUFCMLOADDATA_OUT[7]);
buf B_APUFCMLOADDATA8 (APUFCMLOADDATA[8], APUFCMLOADDATA_OUT[8]);
buf B_APUFCMLOADDATA9 (APUFCMLOADDATA[9], APUFCMLOADDATA_OUT[9]);
buf B_APUFCMLOADDATA10 (APUFCMLOADDATA[10], APUFCMLOADDATA_OUT[10]);
buf B_APUFCMLOADDATA11 (APUFCMLOADDATA[11], APUFCMLOADDATA_OUT[11]);
buf B_APUFCMLOADDATA12 (APUFCMLOADDATA[12], APUFCMLOADDATA_OUT[12]);
buf B_APUFCMLOADDATA13 (APUFCMLOADDATA[13], APUFCMLOADDATA_OUT[13]);
buf B_APUFCMLOADDATA14 (APUFCMLOADDATA[14], APUFCMLOADDATA_OUT[14]);
buf B_APUFCMLOADDATA15 (APUFCMLOADDATA[15], APUFCMLOADDATA_OUT[15]);
buf B_APUFCMLOADDATA16 (APUFCMLOADDATA[16], APUFCMLOADDATA_OUT[16]);
buf B_APUFCMLOADDATA17 (APUFCMLOADDATA[17], APUFCMLOADDATA_OUT[17]);
buf B_APUFCMLOADDATA18 (APUFCMLOADDATA[18], APUFCMLOADDATA_OUT[18]);
buf B_APUFCMLOADDATA19 (APUFCMLOADDATA[19], APUFCMLOADDATA_OUT[19]);
buf B_APUFCMLOADDATA20 (APUFCMLOADDATA[20], APUFCMLOADDATA_OUT[20]);
buf B_APUFCMLOADDATA21 (APUFCMLOADDATA[21], APUFCMLOADDATA_OUT[21]);
buf B_APUFCMLOADDATA22 (APUFCMLOADDATA[22], APUFCMLOADDATA_OUT[22]);
buf B_APUFCMLOADDATA23 (APUFCMLOADDATA[23], APUFCMLOADDATA_OUT[23]);
buf B_APUFCMLOADDATA24 (APUFCMLOADDATA[24], APUFCMLOADDATA_OUT[24]);
buf B_APUFCMLOADDATA25 (APUFCMLOADDATA[25], APUFCMLOADDATA_OUT[25]);
buf B_APUFCMLOADDATA26 (APUFCMLOADDATA[26], APUFCMLOADDATA_OUT[26]);
buf B_APUFCMLOADDATA27 (APUFCMLOADDATA[27], APUFCMLOADDATA_OUT[27]);
buf B_APUFCMLOADDATA28 (APUFCMLOADDATA[28], APUFCMLOADDATA_OUT[28]);
buf B_APUFCMLOADDATA29 (APUFCMLOADDATA[29], APUFCMLOADDATA_OUT[29]);
buf B_APUFCMLOADDATA30 (APUFCMLOADDATA[30], APUFCMLOADDATA_OUT[30]);
buf B_APUFCMLOADDATA31 (APUFCMLOADDATA[31], APUFCMLOADDATA_OUT[31]);
buf B_APUFCMLOADDATA32 (APUFCMLOADDATA[32], APUFCMLOADDATA_OUT[32]);
buf B_APUFCMLOADDATA33 (APUFCMLOADDATA[33], APUFCMLOADDATA_OUT[33]);
buf B_APUFCMLOADDATA34 (APUFCMLOADDATA[34], APUFCMLOADDATA_OUT[34]);
buf B_APUFCMLOADDATA35 (APUFCMLOADDATA[35], APUFCMLOADDATA_OUT[35]);
buf B_APUFCMLOADDATA36 (APUFCMLOADDATA[36], APUFCMLOADDATA_OUT[36]);
buf B_APUFCMLOADDATA37 (APUFCMLOADDATA[37], APUFCMLOADDATA_OUT[37]);
buf B_APUFCMLOADDATA38 (APUFCMLOADDATA[38], APUFCMLOADDATA_OUT[38]);
buf B_APUFCMLOADDATA39 (APUFCMLOADDATA[39], APUFCMLOADDATA_OUT[39]);
buf B_APUFCMLOADDATA40 (APUFCMLOADDATA[40], APUFCMLOADDATA_OUT[40]);
buf B_APUFCMLOADDATA41 (APUFCMLOADDATA[41], APUFCMLOADDATA_OUT[41]);
buf B_APUFCMLOADDATA42 (APUFCMLOADDATA[42], APUFCMLOADDATA_OUT[42]);
buf B_APUFCMLOADDATA43 (APUFCMLOADDATA[43], APUFCMLOADDATA_OUT[43]);
buf B_APUFCMLOADDATA44 (APUFCMLOADDATA[44], APUFCMLOADDATA_OUT[44]);
buf B_APUFCMLOADDATA45 (APUFCMLOADDATA[45], APUFCMLOADDATA_OUT[45]);
buf B_APUFCMLOADDATA46 (APUFCMLOADDATA[46], APUFCMLOADDATA_OUT[46]);
buf B_APUFCMLOADDATA47 (APUFCMLOADDATA[47], APUFCMLOADDATA_OUT[47]);
buf B_APUFCMLOADDATA48 (APUFCMLOADDATA[48], APUFCMLOADDATA_OUT[48]);
buf B_APUFCMLOADDATA49 (APUFCMLOADDATA[49], APUFCMLOADDATA_OUT[49]);
buf B_APUFCMLOADDATA50 (APUFCMLOADDATA[50], APUFCMLOADDATA_OUT[50]);
buf B_APUFCMLOADDATA51 (APUFCMLOADDATA[51], APUFCMLOADDATA_OUT[51]);
buf B_APUFCMLOADDATA52 (APUFCMLOADDATA[52], APUFCMLOADDATA_OUT[52]);
buf B_APUFCMLOADDATA53 (APUFCMLOADDATA[53], APUFCMLOADDATA_OUT[53]);
buf B_APUFCMLOADDATA54 (APUFCMLOADDATA[54], APUFCMLOADDATA_OUT[54]);
buf B_APUFCMLOADDATA55 (APUFCMLOADDATA[55], APUFCMLOADDATA_OUT[55]);
buf B_APUFCMLOADDATA56 (APUFCMLOADDATA[56], APUFCMLOADDATA_OUT[56]);
buf B_APUFCMLOADDATA57 (APUFCMLOADDATA[57], APUFCMLOADDATA_OUT[57]);
buf B_APUFCMLOADDATA58 (APUFCMLOADDATA[58], APUFCMLOADDATA_OUT[58]);
buf B_APUFCMLOADDATA59 (APUFCMLOADDATA[59], APUFCMLOADDATA_OUT[59]);
buf B_APUFCMLOADDATA60 (APUFCMLOADDATA[60], APUFCMLOADDATA_OUT[60]);
buf B_APUFCMLOADDATA61 (APUFCMLOADDATA[61], APUFCMLOADDATA_OUT[61]);
buf B_APUFCMLOADDATA62 (APUFCMLOADDATA[62], APUFCMLOADDATA_OUT[62]);
buf B_APUFCMLOADDATA63 (APUFCMLOADDATA[63], APUFCMLOADDATA_OUT[63]);
buf B_APUFCMLOADDATA64 (APUFCMLOADDATA[64], APUFCMLOADDATA_OUT[64]);
buf B_APUFCMLOADDATA65 (APUFCMLOADDATA[65], APUFCMLOADDATA_OUT[65]);
buf B_APUFCMLOADDATA66 (APUFCMLOADDATA[66], APUFCMLOADDATA_OUT[66]);
buf B_APUFCMLOADDATA67 (APUFCMLOADDATA[67], APUFCMLOADDATA_OUT[67]);
buf B_APUFCMLOADDATA68 (APUFCMLOADDATA[68], APUFCMLOADDATA_OUT[68]);
buf B_APUFCMLOADDATA69 (APUFCMLOADDATA[69], APUFCMLOADDATA_OUT[69]);
buf B_APUFCMLOADDATA70 (APUFCMLOADDATA[70], APUFCMLOADDATA_OUT[70]);
buf B_APUFCMLOADDATA71 (APUFCMLOADDATA[71], APUFCMLOADDATA_OUT[71]);
buf B_APUFCMLOADDATA72 (APUFCMLOADDATA[72], APUFCMLOADDATA_OUT[72]);
buf B_APUFCMLOADDATA73 (APUFCMLOADDATA[73], APUFCMLOADDATA_OUT[73]);
buf B_APUFCMLOADDATA74 (APUFCMLOADDATA[74], APUFCMLOADDATA_OUT[74]);
buf B_APUFCMLOADDATA75 (APUFCMLOADDATA[75], APUFCMLOADDATA_OUT[75]);
buf B_APUFCMLOADDATA76 (APUFCMLOADDATA[76], APUFCMLOADDATA_OUT[76]);
buf B_APUFCMLOADDATA77 (APUFCMLOADDATA[77], APUFCMLOADDATA_OUT[77]);
buf B_APUFCMLOADDATA78 (APUFCMLOADDATA[78], APUFCMLOADDATA_OUT[78]);
buf B_APUFCMLOADDATA79 (APUFCMLOADDATA[79], APUFCMLOADDATA_OUT[79]);
buf B_APUFCMLOADDATA80 (APUFCMLOADDATA[80], APUFCMLOADDATA_OUT[80]);
buf B_APUFCMLOADDATA81 (APUFCMLOADDATA[81], APUFCMLOADDATA_OUT[81]);
buf B_APUFCMLOADDATA82 (APUFCMLOADDATA[82], APUFCMLOADDATA_OUT[82]);
buf B_APUFCMLOADDATA83 (APUFCMLOADDATA[83], APUFCMLOADDATA_OUT[83]);
buf B_APUFCMLOADDATA84 (APUFCMLOADDATA[84], APUFCMLOADDATA_OUT[84]);
buf B_APUFCMLOADDATA85 (APUFCMLOADDATA[85], APUFCMLOADDATA_OUT[85]);
buf B_APUFCMLOADDATA86 (APUFCMLOADDATA[86], APUFCMLOADDATA_OUT[86]);
buf B_APUFCMLOADDATA87 (APUFCMLOADDATA[87], APUFCMLOADDATA_OUT[87]);
buf B_APUFCMLOADDATA88 (APUFCMLOADDATA[88], APUFCMLOADDATA_OUT[88]);
buf B_APUFCMLOADDATA89 (APUFCMLOADDATA[89], APUFCMLOADDATA_OUT[89]);
buf B_APUFCMLOADDATA90 (APUFCMLOADDATA[90], APUFCMLOADDATA_OUT[90]);
buf B_APUFCMLOADDATA91 (APUFCMLOADDATA[91], APUFCMLOADDATA_OUT[91]);
buf B_APUFCMLOADDATA92 (APUFCMLOADDATA[92], APUFCMLOADDATA_OUT[92]);
buf B_APUFCMLOADDATA93 (APUFCMLOADDATA[93], APUFCMLOADDATA_OUT[93]);
buf B_APUFCMLOADDATA94 (APUFCMLOADDATA[94], APUFCMLOADDATA_OUT[94]);
buf B_APUFCMLOADDATA95 (APUFCMLOADDATA[95], APUFCMLOADDATA_OUT[95]);
buf B_APUFCMLOADDATA96 (APUFCMLOADDATA[96], APUFCMLOADDATA_OUT[96]);
buf B_APUFCMLOADDATA97 (APUFCMLOADDATA[97], APUFCMLOADDATA_OUT[97]);
buf B_APUFCMLOADDATA98 (APUFCMLOADDATA[98], APUFCMLOADDATA_OUT[98]);
buf B_APUFCMLOADDATA99 (APUFCMLOADDATA[99], APUFCMLOADDATA_OUT[99]);
buf B_APUFCMLOADDATA100 (APUFCMLOADDATA[100], APUFCMLOADDATA_OUT[100]);
buf B_APUFCMLOADDATA101 (APUFCMLOADDATA[101], APUFCMLOADDATA_OUT[101]);
buf B_APUFCMLOADDATA102 (APUFCMLOADDATA[102], APUFCMLOADDATA_OUT[102]);
buf B_APUFCMLOADDATA103 (APUFCMLOADDATA[103], APUFCMLOADDATA_OUT[103]);
buf B_APUFCMLOADDATA104 (APUFCMLOADDATA[104], APUFCMLOADDATA_OUT[104]);
buf B_APUFCMLOADDATA105 (APUFCMLOADDATA[105], APUFCMLOADDATA_OUT[105]);
buf B_APUFCMLOADDATA106 (APUFCMLOADDATA[106], APUFCMLOADDATA_OUT[106]);
buf B_APUFCMLOADDATA107 (APUFCMLOADDATA[107], APUFCMLOADDATA_OUT[107]);
buf B_APUFCMLOADDATA108 (APUFCMLOADDATA[108], APUFCMLOADDATA_OUT[108]);
buf B_APUFCMLOADDATA109 (APUFCMLOADDATA[109], APUFCMLOADDATA_OUT[109]);
buf B_APUFCMLOADDATA110 (APUFCMLOADDATA[110], APUFCMLOADDATA_OUT[110]);
buf B_APUFCMLOADDATA111 (APUFCMLOADDATA[111], APUFCMLOADDATA_OUT[111]);
buf B_APUFCMLOADDATA112 (APUFCMLOADDATA[112], APUFCMLOADDATA_OUT[112]);
buf B_APUFCMLOADDATA113 (APUFCMLOADDATA[113], APUFCMLOADDATA_OUT[113]);
buf B_APUFCMLOADDATA114 (APUFCMLOADDATA[114], APUFCMLOADDATA_OUT[114]);
buf B_APUFCMLOADDATA115 (APUFCMLOADDATA[115], APUFCMLOADDATA_OUT[115]);
buf B_APUFCMLOADDATA116 (APUFCMLOADDATA[116], APUFCMLOADDATA_OUT[116]);
buf B_APUFCMLOADDATA117 (APUFCMLOADDATA[117], APUFCMLOADDATA_OUT[117]);
buf B_APUFCMLOADDATA118 (APUFCMLOADDATA[118], APUFCMLOADDATA_OUT[118]);
buf B_APUFCMLOADDATA119 (APUFCMLOADDATA[119], APUFCMLOADDATA_OUT[119]);
buf B_APUFCMLOADDATA120 (APUFCMLOADDATA[120], APUFCMLOADDATA_OUT[120]);
buf B_APUFCMLOADDATA121 (APUFCMLOADDATA[121], APUFCMLOADDATA_OUT[121]);
buf B_APUFCMLOADDATA122 (APUFCMLOADDATA[122], APUFCMLOADDATA_OUT[122]);
buf B_APUFCMLOADDATA123 (APUFCMLOADDATA[123], APUFCMLOADDATA_OUT[123]);
buf B_APUFCMLOADDATA124 (APUFCMLOADDATA[124], APUFCMLOADDATA_OUT[124]);
buf B_APUFCMLOADDATA125 (APUFCMLOADDATA[125], APUFCMLOADDATA_OUT[125]);
buf B_APUFCMLOADDATA126 (APUFCMLOADDATA[126], APUFCMLOADDATA_OUT[126]);
buf B_APUFCMLOADDATA127 (APUFCMLOADDATA[127], APUFCMLOADDATA_OUT[127]);
buf B_APUFCMLOADDVALID (APUFCMLOADDVALID, APUFCMLOADDVALID_OUT);
buf B_APUFCMMSRFE0 (APUFCMMSRFE0, APUFCMMSRFE0_OUT);
buf B_APUFCMMSRFE1 (APUFCMMSRFE1, APUFCMMSRFE1_OUT);
buf B_APUFCMNEXTINSTRREADY (APUFCMNEXTINSTRREADY, APUFCMNEXTINSTRREADY_OUT);
buf B_APUFCMOPERANDVALID (APUFCMOPERANDVALID, APUFCMOPERANDVALID_OUT);
buf B_APUFCMRADATA0 (APUFCMRADATA[0], APUFCMRADATA_OUT[0]);
buf B_APUFCMRADATA1 (APUFCMRADATA[1], APUFCMRADATA_OUT[1]);
buf B_APUFCMRADATA2 (APUFCMRADATA[2], APUFCMRADATA_OUT[2]);
buf B_APUFCMRADATA3 (APUFCMRADATA[3], APUFCMRADATA_OUT[3]);
buf B_APUFCMRADATA4 (APUFCMRADATA[4], APUFCMRADATA_OUT[4]);
buf B_APUFCMRADATA5 (APUFCMRADATA[5], APUFCMRADATA_OUT[5]);
buf B_APUFCMRADATA6 (APUFCMRADATA[6], APUFCMRADATA_OUT[6]);
buf B_APUFCMRADATA7 (APUFCMRADATA[7], APUFCMRADATA_OUT[7]);
buf B_APUFCMRADATA8 (APUFCMRADATA[8], APUFCMRADATA_OUT[8]);
buf B_APUFCMRADATA9 (APUFCMRADATA[9], APUFCMRADATA_OUT[9]);
buf B_APUFCMRADATA10 (APUFCMRADATA[10], APUFCMRADATA_OUT[10]);
buf B_APUFCMRADATA11 (APUFCMRADATA[11], APUFCMRADATA_OUT[11]);
buf B_APUFCMRADATA12 (APUFCMRADATA[12], APUFCMRADATA_OUT[12]);
buf B_APUFCMRADATA13 (APUFCMRADATA[13], APUFCMRADATA_OUT[13]);
buf B_APUFCMRADATA14 (APUFCMRADATA[14], APUFCMRADATA_OUT[14]);
buf B_APUFCMRADATA15 (APUFCMRADATA[15], APUFCMRADATA_OUT[15]);
buf B_APUFCMRADATA16 (APUFCMRADATA[16], APUFCMRADATA_OUT[16]);
buf B_APUFCMRADATA17 (APUFCMRADATA[17], APUFCMRADATA_OUT[17]);
buf B_APUFCMRADATA18 (APUFCMRADATA[18], APUFCMRADATA_OUT[18]);
buf B_APUFCMRADATA19 (APUFCMRADATA[19], APUFCMRADATA_OUT[19]);
buf B_APUFCMRADATA20 (APUFCMRADATA[20], APUFCMRADATA_OUT[20]);
buf B_APUFCMRADATA21 (APUFCMRADATA[21], APUFCMRADATA_OUT[21]);
buf B_APUFCMRADATA22 (APUFCMRADATA[22], APUFCMRADATA_OUT[22]);
buf B_APUFCMRADATA23 (APUFCMRADATA[23], APUFCMRADATA_OUT[23]);
buf B_APUFCMRADATA24 (APUFCMRADATA[24], APUFCMRADATA_OUT[24]);
buf B_APUFCMRADATA25 (APUFCMRADATA[25], APUFCMRADATA_OUT[25]);
buf B_APUFCMRADATA26 (APUFCMRADATA[26], APUFCMRADATA_OUT[26]);
buf B_APUFCMRADATA27 (APUFCMRADATA[27], APUFCMRADATA_OUT[27]);
buf B_APUFCMRADATA28 (APUFCMRADATA[28], APUFCMRADATA_OUT[28]);
buf B_APUFCMRADATA29 (APUFCMRADATA[29], APUFCMRADATA_OUT[29]);
buf B_APUFCMRADATA30 (APUFCMRADATA[30], APUFCMRADATA_OUT[30]);
buf B_APUFCMRADATA31 (APUFCMRADATA[31], APUFCMRADATA_OUT[31]);
buf B_APUFCMRBDATA0 (APUFCMRBDATA[0], APUFCMRBDATA_OUT[0]);
buf B_APUFCMRBDATA1 (APUFCMRBDATA[1], APUFCMRBDATA_OUT[1]);
buf B_APUFCMRBDATA2 (APUFCMRBDATA[2], APUFCMRBDATA_OUT[2]);
buf B_APUFCMRBDATA3 (APUFCMRBDATA[3], APUFCMRBDATA_OUT[3]);
buf B_APUFCMRBDATA4 (APUFCMRBDATA[4], APUFCMRBDATA_OUT[4]);
buf B_APUFCMRBDATA5 (APUFCMRBDATA[5], APUFCMRBDATA_OUT[5]);
buf B_APUFCMRBDATA6 (APUFCMRBDATA[6], APUFCMRBDATA_OUT[6]);
buf B_APUFCMRBDATA7 (APUFCMRBDATA[7], APUFCMRBDATA_OUT[7]);
buf B_APUFCMRBDATA8 (APUFCMRBDATA[8], APUFCMRBDATA_OUT[8]);
buf B_APUFCMRBDATA9 (APUFCMRBDATA[9], APUFCMRBDATA_OUT[9]);
buf B_APUFCMRBDATA10 (APUFCMRBDATA[10], APUFCMRBDATA_OUT[10]);
buf B_APUFCMRBDATA11 (APUFCMRBDATA[11], APUFCMRBDATA_OUT[11]);
buf B_APUFCMRBDATA12 (APUFCMRBDATA[12], APUFCMRBDATA_OUT[12]);
buf B_APUFCMRBDATA13 (APUFCMRBDATA[13], APUFCMRBDATA_OUT[13]);
buf B_APUFCMRBDATA14 (APUFCMRBDATA[14], APUFCMRBDATA_OUT[14]);
buf B_APUFCMRBDATA15 (APUFCMRBDATA[15], APUFCMRBDATA_OUT[15]);
buf B_APUFCMRBDATA16 (APUFCMRBDATA[16], APUFCMRBDATA_OUT[16]);
buf B_APUFCMRBDATA17 (APUFCMRBDATA[17], APUFCMRBDATA_OUT[17]);
buf B_APUFCMRBDATA18 (APUFCMRBDATA[18], APUFCMRBDATA_OUT[18]);
buf B_APUFCMRBDATA19 (APUFCMRBDATA[19], APUFCMRBDATA_OUT[19]);
buf B_APUFCMRBDATA20 (APUFCMRBDATA[20], APUFCMRBDATA_OUT[20]);
buf B_APUFCMRBDATA21 (APUFCMRBDATA[21], APUFCMRBDATA_OUT[21]);
buf B_APUFCMRBDATA22 (APUFCMRBDATA[22], APUFCMRBDATA_OUT[22]);
buf B_APUFCMRBDATA23 (APUFCMRBDATA[23], APUFCMRBDATA_OUT[23]);
buf B_APUFCMRBDATA24 (APUFCMRBDATA[24], APUFCMRBDATA_OUT[24]);
buf B_APUFCMRBDATA25 (APUFCMRBDATA[25], APUFCMRBDATA_OUT[25]);
buf B_APUFCMRBDATA26 (APUFCMRBDATA[26], APUFCMRBDATA_OUT[26]);
buf B_APUFCMRBDATA27 (APUFCMRBDATA[27], APUFCMRBDATA_OUT[27]);
buf B_APUFCMRBDATA28 (APUFCMRBDATA[28], APUFCMRBDATA_OUT[28]);
buf B_APUFCMRBDATA29 (APUFCMRBDATA[29], APUFCMRBDATA_OUT[29]);
buf B_APUFCMRBDATA30 (APUFCMRBDATA[30], APUFCMRBDATA_OUT[30]);
buf B_APUFCMRBDATA31 (APUFCMRBDATA[31], APUFCMRBDATA_OUT[31]);
buf B_APUFCMWRITEBACKOK (APUFCMWRITEBACKOK, APUFCMWRITEBACKOK_OUT);
buf B_C440CPMCORESLEEPREQ (C440CPMCORESLEEPREQ, C440CPMCORESLEEPREQ_OUT);
buf B_C440CPMDECIRPTREQ (C440CPMDECIRPTREQ, C440CPMDECIRPTREQ_OUT);
buf B_C440CPMFITIRPTREQ (C440CPMFITIRPTREQ, C440CPMFITIRPTREQ_OUT);
buf B_C440CPMMSRCE (C440CPMMSRCE, C440CPMMSRCE_OUT);
buf B_C440CPMMSREE (C440CPMMSREE, C440CPMMSREE_OUT);
buf B_C440CPMTIMERRESETREQ (C440CPMTIMERRESETREQ, C440CPMTIMERRESETREQ_OUT);
buf B_C440CPMWDIRPTREQ (C440CPMWDIRPTREQ, C440CPMWDIRPTREQ_OUT);
buf B_C440DBGSYSTEMCONTROL0 (C440DBGSYSTEMCONTROL[0], C440DBGSYSTEMCONTROL_OUT[0]);
buf B_C440DBGSYSTEMCONTROL1 (C440DBGSYSTEMCONTROL[1], C440DBGSYSTEMCONTROL_OUT[1]);
buf B_C440DBGSYSTEMCONTROL2 (C440DBGSYSTEMCONTROL[2], C440DBGSYSTEMCONTROL_OUT[2]);
buf B_C440DBGSYSTEMCONTROL3 (C440DBGSYSTEMCONTROL[3], C440DBGSYSTEMCONTROL_OUT[3]);
buf B_C440DBGSYSTEMCONTROL4 (C440DBGSYSTEMCONTROL[4], C440DBGSYSTEMCONTROL_OUT[4]);
buf B_C440DBGSYSTEMCONTROL5 (C440DBGSYSTEMCONTROL[5], C440DBGSYSTEMCONTROL_OUT[5]);
buf B_C440DBGSYSTEMCONTROL6 (C440DBGSYSTEMCONTROL[6], C440DBGSYSTEMCONTROL_OUT[6]);
buf B_C440DBGSYSTEMCONTROL7 (C440DBGSYSTEMCONTROL[7], C440DBGSYSTEMCONTROL_OUT[7]);
buf B_C440JTGTDO (C440JTGTDO, C440JTGTDO_OUT);
buf B_C440JTGTDOEN (C440JTGTDOEN, C440JTGTDOEN_OUT);
buf B_C440MACHINECHECK (C440MACHINECHECK, C440MACHINECHECK_OUT);
buf B_C440RSTCHIPRESETREQ (C440RSTCHIPRESETREQ, C440RSTCHIPRESETREQ_OUT);
buf B_C440RSTCORERESETREQ (C440RSTCORERESETREQ, C440RSTCORERESETREQ_OUT);
buf B_C440RSTSYSTEMRESETREQ (C440RSTSYSTEMRESETREQ, C440RSTSYSTEMRESETREQ_OUT);
buf B_C440TRCBRANCHSTATUS0 (C440TRCBRANCHSTATUS[0], C440TRCBRANCHSTATUS_OUT[0]);
buf B_C440TRCBRANCHSTATUS1 (C440TRCBRANCHSTATUS[1], C440TRCBRANCHSTATUS_OUT[1]);
buf B_C440TRCBRANCHSTATUS2 (C440TRCBRANCHSTATUS[2], C440TRCBRANCHSTATUS_OUT[2]);
buf B_C440TRCCYCLE (C440TRCCYCLE, C440TRCCYCLE_OUT);
buf B_C440TRCEXECUTIONSTATUS0 (C440TRCEXECUTIONSTATUS[0], C440TRCEXECUTIONSTATUS_OUT[0]);
buf B_C440TRCEXECUTIONSTATUS1 (C440TRCEXECUTIONSTATUS[1], C440TRCEXECUTIONSTATUS_OUT[1]);
buf B_C440TRCEXECUTIONSTATUS2 (C440TRCEXECUTIONSTATUS[2], C440TRCEXECUTIONSTATUS_OUT[2]);
buf B_C440TRCEXECUTIONSTATUS3 (C440TRCEXECUTIONSTATUS[3], C440TRCEXECUTIONSTATUS_OUT[3]);
buf B_C440TRCEXECUTIONSTATUS4 (C440TRCEXECUTIONSTATUS[4], C440TRCEXECUTIONSTATUS_OUT[4]);
buf B_C440TRCTRACESTATUS0 (C440TRCTRACESTATUS[0], C440TRCTRACESTATUS_OUT[0]);
buf B_C440TRCTRACESTATUS1 (C440TRCTRACESTATUS[1], C440TRCTRACESTATUS_OUT[1]);
buf B_C440TRCTRACESTATUS2 (C440TRCTRACESTATUS[2], C440TRCTRACESTATUS_OUT[2]);
buf B_C440TRCTRACESTATUS3 (C440TRCTRACESTATUS[3], C440TRCTRACESTATUS_OUT[3]);
buf B_C440TRCTRACESTATUS4 (C440TRCTRACESTATUS[4], C440TRCTRACESTATUS_OUT[4]);
buf B_C440TRCTRACESTATUS5 (C440TRCTRACESTATUS[5], C440TRCTRACESTATUS_OUT[5]);
buf B_C440TRCTRACESTATUS6 (C440TRCTRACESTATUS[6], C440TRCTRACESTATUS_OUT[6]);
buf B_C440TRCTRIGGEREVENTOUT (C440TRCTRIGGEREVENTOUT, C440TRCTRIGGEREVENTOUT_OUT);
buf B_C440TRCTRIGGEREVENTTYPE0 (C440TRCTRIGGEREVENTTYPE[0], C440TRCTRIGGEREVENTTYPE_OUT[0]);
buf B_C440TRCTRIGGEREVENTTYPE1 (C440TRCTRIGGEREVENTTYPE[1], C440TRCTRIGGEREVENTTYPE_OUT[1]);
buf B_C440TRCTRIGGEREVENTTYPE2 (C440TRCTRIGGEREVENTTYPE[2], C440TRCTRIGGEREVENTTYPE_OUT[2]);
buf B_C440TRCTRIGGEREVENTTYPE3 (C440TRCTRIGGEREVENTTYPE[3], C440TRCTRIGGEREVENTTYPE_OUT[3]);
buf B_C440TRCTRIGGEREVENTTYPE4 (C440TRCTRIGGEREVENTTYPE[4], C440TRCTRIGGEREVENTTYPE_OUT[4]);
buf B_C440TRCTRIGGEREVENTTYPE5 (C440TRCTRIGGEREVENTTYPE[5], C440TRCTRIGGEREVENTTYPE_OUT[5]);
buf B_C440TRCTRIGGEREVENTTYPE6 (C440TRCTRIGGEREVENTTYPE[6], C440TRCTRIGGEREVENTTYPE_OUT[6]);
buf B_C440TRCTRIGGEREVENTTYPE7 (C440TRCTRIGGEREVENTTYPE[7], C440TRCTRIGGEREVENTTYPE_OUT[7]);
buf B_C440TRCTRIGGEREVENTTYPE8 (C440TRCTRIGGEREVENTTYPE[8], C440TRCTRIGGEREVENTTYPE_OUT[8]);
buf B_C440TRCTRIGGEREVENTTYPE9 (C440TRCTRIGGEREVENTTYPE[9], C440TRCTRIGGEREVENTTYPE_OUT[9]);
buf B_C440TRCTRIGGEREVENTTYPE10 (C440TRCTRIGGEREVENTTYPE[10], C440TRCTRIGGEREVENTTYPE_OUT[10]);
buf B_C440TRCTRIGGEREVENTTYPE11 (C440TRCTRIGGEREVENTTYPE[11], C440TRCTRIGGEREVENTTYPE_OUT[11]);
buf B_C440TRCTRIGGEREVENTTYPE12 (C440TRCTRIGGEREVENTTYPE[12], C440TRCTRIGGEREVENTTYPE_OUT[12]);
buf B_C440TRCTRIGGEREVENTTYPE13 (C440TRCTRIGGEREVENTTYPE[13], C440TRCTRIGGEREVENTTYPE_OUT[13]);
buf B_MIMCADDRESS0 (MIMCADDRESS[0], MIMCADDRESS_OUT[0]);
buf B_MIMCADDRESS1 (MIMCADDRESS[1], MIMCADDRESS_OUT[1]);
buf B_MIMCADDRESS2 (MIMCADDRESS[2], MIMCADDRESS_OUT[2]);
buf B_MIMCADDRESS3 (MIMCADDRESS[3], MIMCADDRESS_OUT[3]);
buf B_MIMCADDRESS4 (MIMCADDRESS[4], MIMCADDRESS_OUT[4]);
buf B_MIMCADDRESS5 (MIMCADDRESS[5], MIMCADDRESS_OUT[5]);
buf B_MIMCADDRESS6 (MIMCADDRESS[6], MIMCADDRESS_OUT[6]);
buf B_MIMCADDRESS7 (MIMCADDRESS[7], MIMCADDRESS_OUT[7]);
buf B_MIMCADDRESS8 (MIMCADDRESS[8], MIMCADDRESS_OUT[8]);
buf B_MIMCADDRESS9 (MIMCADDRESS[9], MIMCADDRESS_OUT[9]);
buf B_MIMCADDRESS10 (MIMCADDRESS[10], MIMCADDRESS_OUT[10]);
buf B_MIMCADDRESS11 (MIMCADDRESS[11], MIMCADDRESS_OUT[11]);
buf B_MIMCADDRESS12 (MIMCADDRESS[12], MIMCADDRESS_OUT[12]);
buf B_MIMCADDRESS13 (MIMCADDRESS[13], MIMCADDRESS_OUT[13]);
buf B_MIMCADDRESS14 (MIMCADDRESS[14], MIMCADDRESS_OUT[14]);
buf B_MIMCADDRESS15 (MIMCADDRESS[15], MIMCADDRESS_OUT[15]);
buf B_MIMCADDRESS16 (MIMCADDRESS[16], MIMCADDRESS_OUT[16]);
buf B_MIMCADDRESS17 (MIMCADDRESS[17], MIMCADDRESS_OUT[17]);
buf B_MIMCADDRESS18 (MIMCADDRESS[18], MIMCADDRESS_OUT[18]);
buf B_MIMCADDRESS19 (MIMCADDRESS[19], MIMCADDRESS_OUT[19]);
buf B_MIMCADDRESS20 (MIMCADDRESS[20], MIMCADDRESS_OUT[20]);
buf B_MIMCADDRESS21 (MIMCADDRESS[21], MIMCADDRESS_OUT[21]);
buf B_MIMCADDRESS22 (MIMCADDRESS[22], MIMCADDRESS_OUT[22]);
buf B_MIMCADDRESS23 (MIMCADDRESS[23], MIMCADDRESS_OUT[23]);
buf B_MIMCADDRESS24 (MIMCADDRESS[24], MIMCADDRESS_OUT[24]);
buf B_MIMCADDRESS25 (MIMCADDRESS[25], MIMCADDRESS_OUT[25]);
buf B_MIMCADDRESS26 (MIMCADDRESS[26], MIMCADDRESS_OUT[26]);
buf B_MIMCADDRESS27 (MIMCADDRESS[27], MIMCADDRESS_OUT[27]);
buf B_MIMCADDRESS28 (MIMCADDRESS[28], MIMCADDRESS_OUT[28]);
buf B_MIMCADDRESS29 (MIMCADDRESS[29], MIMCADDRESS_OUT[29]);
buf B_MIMCADDRESS30 (MIMCADDRESS[30], MIMCADDRESS_OUT[30]);
buf B_MIMCADDRESS31 (MIMCADDRESS[31], MIMCADDRESS_OUT[31]);
buf B_MIMCADDRESS32 (MIMCADDRESS[32], MIMCADDRESS_OUT[32]);
buf B_MIMCADDRESS33 (MIMCADDRESS[33], MIMCADDRESS_OUT[33]);
buf B_MIMCADDRESS34 (MIMCADDRESS[34], MIMCADDRESS_OUT[34]);
buf B_MIMCADDRESS35 (MIMCADDRESS[35], MIMCADDRESS_OUT[35]);
buf B_MIMCADDRESSVALID (MIMCADDRESSVALID, MIMCADDRESSVALID_OUT);
buf B_MIMCBANKCONFLICT (MIMCBANKCONFLICT, MIMCBANKCONFLICT_OUT);
buf B_MIMCBYTEENABLE0 (MIMCBYTEENABLE[0], MIMCBYTEENABLE_OUT[0]);
buf B_MIMCBYTEENABLE1 (MIMCBYTEENABLE[1], MIMCBYTEENABLE_OUT[1]);
buf B_MIMCBYTEENABLE2 (MIMCBYTEENABLE[2], MIMCBYTEENABLE_OUT[2]);
buf B_MIMCBYTEENABLE3 (MIMCBYTEENABLE[3], MIMCBYTEENABLE_OUT[3]);
buf B_MIMCBYTEENABLE4 (MIMCBYTEENABLE[4], MIMCBYTEENABLE_OUT[4]);
buf B_MIMCBYTEENABLE5 (MIMCBYTEENABLE[5], MIMCBYTEENABLE_OUT[5]);
buf B_MIMCBYTEENABLE6 (MIMCBYTEENABLE[6], MIMCBYTEENABLE_OUT[6]);
buf B_MIMCBYTEENABLE7 (MIMCBYTEENABLE[7], MIMCBYTEENABLE_OUT[7]);
buf B_MIMCBYTEENABLE8 (MIMCBYTEENABLE[8], MIMCBYTEENABLE_OUT[8]);
buf B_MIMCBYTEENABLE9 (MIMCBYTEENABLE[9], MIMCBYTEENABLE_OUT[9]);
buf B_MIMCBYTEENABLE10 (MIMCBYTEENABLE[10], MIMCBYTEENABLE_OUT[10]);
buf B_MIMCBYTEENABLE11 (MIMCBYTEENABLE[11], MIMCBYTEENABLE_OUT[11]);
buf B_MIMCBYTEENABLE12 (MIMCBYTEENABLE[12], MIMCBYTEENABLE_OUT[12]);
buf B_MIMCBYTEENABLE13 (MIMCBYTEENABLE[13], MIMCBYTEENABLE_OUT[13]);
buf B_MIMCBYTEENABLE14 (MIMCBYTEENABLE[14], MIMCBYTEENABLE_OUT[14]);
buf B_MIMCBYTEENABLE15 (MIMCBYTEENABLE[15], MIMCBYTEENABLE_OUT[15]);
buf B_MIMCREADNOTWRITE (MIMCREADNOTWRITE, MIMCREADNOTWRITE_OUT);
buf B_MIMCROWCONFLICT (MIMCROWCONFLICT, MIMCROWCONFLICT_OUT);
buf B_MIMCWRITEDATA0 (MIMCWRITEDATA[0], MIMCWRITEDATA_OUT[0]);
buf B_MIMCWRITEDATA1 (MIMCWRITEDATA[1], MIMCWRITEDATA_OUT[1]);
buf B_MIMCWRITEDATA2 (MIMCWRITEDATA[2], MIMCWRITEDATA_OUT[2]);
buf B_MIMCWRITEDATA3 (MIMCWRITEDATA[3], MIMCWRITEDATA_OUT[3]);
buf B_MIMCWRITEDATA4 (MIMCWRITEDATA[4], MIMCWRITEDATA_OUT[4]);
buf B_MIMCWRITEDATA5 (MIMCWRITEDATA[5], MIMCWRITEDATA_OUT[5]);
buf B_MIMCWRITEDATA6 (MIMCWRITEDATA[6], MIMCWRITEDATA_OUT[6]);
buf B_MIMCWRITEDATA7 (MIMCWRITEDATA[7], MIMCWRITEDATA_OUT[7]);
buf B_MIMCWRITEDATA8 (MIMCWRITEDATA[8], MIMCWRITEDATA_OUT[8]);
buf B_MIMCWRITEDATA9 (MIMCWRITEDATA[9], MIMCWRITEDATA_OUT[9]);
buf B_MIMCWRITEDATA10 (MIMCWRITEDATA[10], MIMCWRITEDATA_OUT[10]);
buf B_MIMCWRITEDATA11 (MIMCWRITEDATA[11], MIMCWRITEDATA_OUT[11]);
buf B_MIMCWRITEDATA12 (MIMCWRITEDATA[12], MIMCWRITEDATA_OUT[12]);
buf B_MIMCWRITEDATA13 (MIMCWRITEDATA[13], MIMCWRITEDATA_OUT[13]);
buf B_MIMCWRITEDATA14 (MIMCWRITEDATA[14], MIMCWRITEDATA_OUT[14]);
buf B_MIMCWRITEDATA15 (MIMCWRITEDATA[15], MIMCWRITEDATA_OUT[15]);
buf B_MIMCWRITEDATA16 (MIMCWRITEDATA[16], MIMCWRITEDATA_OUT[16]);
buf B_MIMCWRITEDATA17 (MIMCWRITEDATA[17], MIMCWRITEDATA_OUT[17]);
buf B_MIMCWRITEDATA18 (MIMCWRITEDATA[18], MIMCWRITEDATA_OUT[18]);
buf B_MIMCWRITEDATA19 (MIMCWRITEDATA[19], MIMCWRITEDATA_OUT[19]);
buf B_MIMCWRITEDATA20 (MIMCWRITEDATA[20], MIMCWRITEDATA_OUT[20]);
buf B_MIMCWRITEDATA21 (MIMCWRITEDATA[21], MIMCWRITEDATA_OUT[21]);
buf B_MIMCWRITEDATA22 (MIMCWRITEDATA[22], MIMCWRITEDATA_OUT[22]);
buf B_MIMCWRITEDATA23 (MIMCWRITEDATA[23], MIMCWRITEDATA_OUT[23]);
buf B_MIMCWRITEDATA24 (MIMCWRITEDATA[24], MIMCWRITEDATA_OUT[24]);
buf B_MIMCWRITEDATA25 (MIMCWRITEDATA[25], MIMCWRITEDATA_OUT[25]);
buf B_MIMCWRITEDATA26 (MIMCWRITEDATA[26], MIMCWRITEDATA_OUT[26]);
buf B_MIMCWRITEDATA27 (MIMCWRITEDATA[27], MIMCWRITEDATA_OUT[27]);
buf B_MIMCWRITEDATA28 (MIMCWRITEDATA[28], MIMCWRITEDATA_OUT[28]);
buf B_MIMCWRITEDATA29 (MIMCWRITEDATA[29], MIMCWRITEDATA_OUT[29]);
buf B_MIMCWRITEDATA30 (MIMCWRITEDATA[30], MIMCWRITEDATA_OUT[30]);
buf B_MIMCWRITEDATA31 (MIMCWRITEDATA[31], MIMCWRITEDATA_OUT[31]);
buf B_MIMCWRITEDATA32 (MIMCWRITEDATA[32], MIMCWRITEDATA_OUT[32]);
buf B_MIMCWRITEDATA33 (MIMCWRITEDATA[33], MIMCWRITEDATA_OUT[33]);
buf B_MIMCWRITEDATA34 (MIMCWRITEDATA[34], MIMCWRITEDATA_OUT[34]);
buf B_MIMCWRITEDATA35 (MIMCWRITEDATA[35], MIMCWRITEDATA_OUT[35]);
buf B_MIMCWRITEDATA36 (MIMCWRITEDATA[36], MIMCWRITEDATA_OUT[36]);
buf B_MIMCWRITEDATA37 (MIMCWRITEDATA[37], MIMCWRITEDATA_OUT[37]);
buf B_MIMCWRITEDATA38 (MIMCWRITEDATA[38], MIMCWRITEDATA_OUT[38]);
buf B_MIMCWRITEDATA39 (MIMCWRITEDATA[39], MIMCWRITEDATA_OUT[39]);
buf B_MIMCWRITEDATA40 (MIMCWRITEDATA[40], MIMCWRITEDATA_OUT[40]);
buf B_MIMCWRITEDATA41 (MIMCWRITEDATA[41], MIMCWRITEDATA_OUT[41]);
buf B_MIMCWRITEDATA42 (MIMCWRITEDATA[42], MIMCWRITEDATA_OUT[42]);
buf B_MIMCWRITEDATA43 (MIMCWRITEDATA[43], MIMCWRITEDATA_OUT[43]);
buf B_MIMCWRITEDATA44 (MIMCWRITEDATA[44], MIMCWRITEDATA_OUT[44]);
buf B_MIMCWRITEDATA45 (MIMCWRITEDATA[45], MIMCWRITEDATA_OUT[45]);
buf B_MIMCWRITEDATA46 (MIMCWRITEDATA[46], MIMCWRITEDATA_OUT[46]);
buf B_MIMCWRITEDATA47 (MIMCWRITEDATA[47], MIMCWRITEDATA_OUT[47]);
buf B_MIMCWRITEDATA48 (MIMCWRITEDATA[48], MIMCWRITEDATA_OUT[48]);
buf B_MIMCWRITEDATA49 (MIMCWRITEDATA[49], MIMCWRITEDATA_OUT[49]);
buf B_MIMCWRITEDATA50 (MIMCWRITEDATA[50], MIMCWRITEDATA_OUT[50]);
buf B_MIMCWRITEDATA51 (MIMCWRITEDATA[51], MIMCWRITEDATA_OUT[51]);
buf B_MIMCWRITEDATA52 (MIMCWRITEDATA[52], MIMCWRITEDATA_OUT[52]);
buf B_MIMCWRITEDATA53 (MIMCWRITEDATA[53], MIMCWRITEDATA_OUT[53]);
buf B_MIMCWRITEDATA54 (MIMCWRITEDATA[54], MIMCWRITEDATA_OUT[54]);
buf B_MIMCWRITEDATA55 (MIMCWRITEDATA[55], MIMCWRITEDATA_OUT[55]);
buf B_MIMCWRITEDATA56 (MIMCWRITEDATA[56], MIMCWRITEDATA_OUT[56]);
buf B_MIMCWRITEDATA57 (MIMCWRITEDATA[57], MIMCWRITEDATA_OUT[57]);
buf B_MIMCWRITEDATA58 (MIMCWRITEDATA[58], MIMCWRITEDATA_OUT[58]);
buf B_MIMCWRITEDATA59 (MIMCWRITEDATA[59], MIMCWRITEDATA_OUT[59]);
buf B_MIMCWRITEDATA60 (MIMCWRITEDATA[60], MIMCWRITEDATA_OUT[60]);
buf B_MIMCWRITEDATA61 (MIMCWRITEDATA[61], MIMCWRITEDATA_OUT[61]);
buf B_MIMCWRITEDATA62 (MIMCWRITEDATA[62], MIMCWRITEDATA_OUT[62]);
buf B_MIMCWRITEDATA63 (MIMCWRITEDATA[63], MIMCWRITEDATA_OUT[63]);
buf B_MIMCWRITEDATA64 (MIMCWRITEDATA[64], MIMCWRITEDATA_OUT[64]);
buf B_MIMCWRITEDATA65 (MIMCWRITEDATA[65], MIMCWRITEDATA_OUT[65]);
buf B_MIMCWRITEDATA66 (MIMCWRITEDATA[66], MIMCWRITEDATA_OUT[66]);
buf B_MIMCWRITEDATA67 (MIMCWRITEDATA[67], MIMCWRITEDATA_OUT[67]);
buf B_MIMCWRITEDATA68 (MIMCWRITEDATA[68], MIMCWRITEDATA_OUT[68]);
buf B_MIMCWRITEDATA69 (MIMCWRITEDATA[69], MIMCWRITEDATA_OUT[69]);
buf B_MIMCWRITEDATA70 (MIMCWRITEDATA[70], MIMCWRITEDATA_OUT[70]);
buf B_MIMCWRITEDATA71 (MIMCWRITEDATA[71], MIMCWRITEDATA_OUT[71]);
buf B_MIMCWRITEDATA72 (MIMCWRITEDATA[72], MIMCWRITEDATA_OUT[72]);
buf B_MIMCWRITEDATA73 (MIMCWRITEDATA[73], MIMCWRITEDATA_OUT[73]);
buf B_MIMCWRITEDATA74 (MIMCWRITEDATA[74], MIMCWRITEDATA_OUT[74]);
buf B_MIMCWRITEDATA75 (MIMCWRITEDATA[75], MIMCWRITEDATA_OUT[75]);
buf B_MIMCWRITEDATA76 (MIMCWRITEDATA[76], MIMCWRITEDATA_OUT[76]);
buf B_MIMCWRITEDATA77 (MIMCWRITEDATA[77], MIMCWRITEDATA_OUT[77]);
buf B_MIMCWRITEDATA78 (MIMCWRITEDATA[78], MIMCWRITEDATA_OUT[78]);
buf B_MIMCWRITEDATA79 (MIMCWRITEDATA[79], MIMCWRITEDATA_OUT[79]);
buf B_MIMCWRITEDATA80 (MIMCWRITEDATA[80], MIMCWRITEDATA_OUT[80]);
buf B_MIMCWRITEDATA81 (MIMCWRITEDATA[81], MIMCWRITEDATA_OUT[81]);
buf B_MIMCWRITEDATA82 (MIMCWRITEDATA[82], MIMCWRITEDATA_OUT[82]);
buf B_MIMCWRITEDATA83 (MIMCWRITEDATA[83], MIMCWRITEDATA_OUT[83]);
buf B_MIMCWRITEDATA84 (MIMCWRITEDATA[84], MIMCWRITEDATA_OUT[84]);
buf B_MIMCWRITEDATA85 (MIMCWRITEDATA[85], MIMCWRITEDATA_OUT[85]);
buf B_MIMCWRITEDATA86 (MIMCWRITEDATA[86], MIMCWRITEDATA_OUT[86]);
buf B_MIMCWRITEDATA87 (MIMCWRITEDATA[87], MIMCWRITEDATA_OUT[87]);
buf B_MIMCWRITEDATA88 (MIMCWRITEDATA[88], MIMCWRITEDATA_OUT[88]);
buf B_MIMCWRITEDATA89 (MIMCWRITEDATA[89], MIMCWRITEDATA_OUT[89]);
buf B_MIMCWRITEDATA90 (MIMCWRITEDATA[90], MIMCWRITEDATA_OUT[90]);
buf B_MIMCWRITEDATA91 (MIMCWRITEDATA[91], MIMCWRITEDATA_OUT[91]);
buf B_MIMCWRITEDATA92 (MIMCWRITEDATA[92], MIMCWRITEDATA_OUT[92]);
buf B_MIMCWRITEDATA93 (MIMCWRITEDATA[93], MIMCWRITEDATA_OUT[93]);
buf B_MIMCWRITEDATA94 (MIMCWRITEDATA[94], MIMCWRITEDATA_OUT[94]);
buf B_MIMCWRITEDATA95 (MIMCWRITEDATA[95], MIMCWRITEDATA_OUT[95]);
buf B_MIMCWRITEDATA96 (MIMCWRITEDATA[96], MIMCWRITEDATA_OUT[96]);
buf B_MIMCWRITEDATA97 (MIMCWRITEDATA[97], MIMCWRITEDATA_OUT[97]);
buf B_MIMCWRITEDATA98 (MIMCWRITEDATA[98], MIMCWRITEDATA_OUT[98]);
buf B_MIMCWRITEDATA99 (MIMCWRITEDATA[99], MIMCWRITEDATA_OUT[99]);
buf B_MIMCWRITEDATA100 (MIMCWRITEDATA[100], MIMCWRITEDATA_OUT[100]);
buf B_MIMCWRITEDATA101 (MIMCWRITEDATA[101], MIMCWRITEDATA_OUT[101]);
buf B_MIMCWRITEDATA102 (MIMCWRITEDATA[102], MIMCWRITEDATA_OUT[102]);
buf B_MIMCWRITEDATA103 (MIMCWRITEDATA[103], MIMCWRITEDATA_OUT[103]);
buf B_MIMCWRITEDATA104 (MIMCWRITEDATA[104], MIMCWRITEDATA_OUT[104]);
buf B_MIMCWRITEDATA105 (MIMCWRITEDATA[105], MIMCWRITEDATA_OUT[105]);
buf B_MIMCWRITEDATA106 (MIMCWRITEDATA[106], MIMCWRITEDATA_OUT[106]);
buf B_MIMCWRITEDATA107 (MIMCWRITEDATA[107], MIMCWRITEDATA_OUT[107]);
buf B_MIMCWRITEDATA108 (MIMCWRITEDATA[108], MIMCWRITEDATA_OUT[108]);
buf B_MIMCWRITEDATA109 (MIMCWRITEDATA[109], MIMCWRITEDATA_OUT[109]);
buf B_MIMCWRITEDATA110 (MIMCWRITEDATA[110], MIMCWRITEDATA_OUT[110]);
buf B_MIMCWRITEDATA111 (MIMCWRITEDATA[111], MIMCWRITEDATA_OUT[111]);
buf B_MIMCWRITEDATA112 (MIMCWRITEDATA[112], MIMCWRITEDATA_OUT[112]);
buf B_MIMCWRITEDATA113 (MIMCWRITEDATA[113], MIMCWRITEDATA_OUT[113]);
buf B_MIMCWRITEDATA114 (MIMCWRITEDATA[114], MIMCWRITEDATA_OUT[114]);
buf B_MIMCWRITEDATA115 (MIMCWRITEDATA[115], MIMCWRITEDATA_OUT[115]);
buf B_MIMCWRITEDATA116 (MIMCWRITEDATA[116], MIMCWRITEDATA_OUT[116]);
buf B_MIMCWRITEDATA117 (MIMCWRITEDATA[117], MIMCWRITEDATA_OUT[117]);
buf B_MIMCWRITEDATA118 (MIMCWRITEDATA[118], MIMCWRITEDATA_OUT[118]);
buf B_MIMCWRITEDATA119 (MIMCWRITEDATA[119], MIMCWRITEDATA_OUT[119]);
buf B_MIMCWRITEDATA120 (MIMCWRITEDATA[120], MIMCWRITEDATA_OUT[120]);
buf B_MIMCWRITEDATA121 (MIMCWRITEDATA[121], MIMCWRITEDATA_OUT[121]);
buf B_MIMCWRITEDATA122 (MIMCWRITEDATA[122], MIMCWRITEDATA_OUT[122]);
buf B_MIMCWRITEDATA123 (MIMCWRITEDATA[123], MIMCWRITEDATA_OUT[123]);
buf B_MIMCWRITEDATA124 (MIMCWRITEDATA[124], MIMCWRITEDATA_OUT[124]);
buf B_MIMCWRITEDATA125 (MIMCWRITEDATA[125], MIMCWRITEDATA_OUT[125]);
buf B_MIMCWRITEDATA126 (MIMCWRITEDATA[126], MIMCWRITEDATA_OUT[126]);
buf B_MIMCWRITEDATA127 (MIMCWRITEDATA[127], MIMCWRITEDATA_OUT[127]);
buf B_MIMCWRITEDATAVALID (MIMCWRITEDATAVALID, MIMCWRITEDATAVALID_OUT);
buf B_PPCCPMINTERCONNECTBUSY (PPCCPMINTERCONNECTBUSY, PPCCPMINTERCONNECTBUSY_OUT);
buf B_PPCDSDCRACK (PPCDSDCRACK, PPCDSDCRACK_OUT);
buf B_PPCDSDCRTIMEOUTWAIT (PPCDSDCRTIMEOUTWAIT, PPCDSDCRTIMEOUTWAIT_OUT);
buf B_PPCDSDCRDBUSIN0 (PPCDSDCRDBUSIN[0], PPCDSDCRDBUSIN_OUT[0]);
buf B_PPCDSDCRDBUSIN1 (PPCDSDCRDBUSIN[1], PPCDSDCRDBUSIN_OUT[1]);
buf B_PPCDSDCRDBUSIN2 (PPCDSDCRDBUSIN[2], PPCDSDCRDBUSIN_OUT[2]);
buf B_PPCDSDCRDBUSIN3 (PPCDSDCRDBUSIN[3], PPCDSDCRDBUSIN_OUT[3]);
buf B_PPCDSDCRDBUSIN4 (PPCDSDCRDBUSIN[4], PPCDSDCRDBUSIN_OUT[4]);
buf B_PPCDSDCRDBUSIN5 (PPCDSDCRDBUSIN[5], PPCDSDCRDBUSIN_OUT[5]);
buf B_PPCDSDCRDBUSIN6 (PPCDSDCRDBUSIN[6], PPCDSDCRDBUSIN_OUT[6]);
buf B_PPCDSDCRDBUSIN7 (PPCDSDCRDBUSIN[7], PPCDSDCRDBUSIN_OUT[7]);
buf B_PPCDSDCRDBUSIN8 (PPCDSDCRDBUSIN[8], PPCDSDCRDBUSIN_OUT[8]);
buf B_PPCDSDCRDBUSIN9 (PPCDSDCRDBUSIN[9], PPCDSDCRDBUSIN_OUT[9]);
buf B_PPCDSDCRDBUSIN10 (PPCDSDCRDBUSIN[10], PPCDSDCRDBUSIN_OUT[10]);
buf B_PPCDSDCRDBUSIN11 (PPCDSDCRDBUSIN[11], PPCDSDCRDBUSIN_OUT[11]);
buf B_PPCDSDCRDBUSIN12 (PPCDSDCRDBUSIN[12], PPCDSDCRDBUSIN_OUT[12]);
buf B_PPCDSDCRDBUSIN13 (PPCDSDCRDBUSIN[13], PPCDSDCRDBUSIN_OUT[13]);
buf B_PPCDSDCRDBUSIN14 (PPCDSDCRDBUSIN[14], PPCDSDCRDBUSIN_OUT[14]);
buf B_PPCDSDCRDBUSIN15 (PPCDSDCRDBUSIN[15], PPCDSDCRDBUSIN_OUT[15]);
buf B_PPCDSDCRDBUSIN16 (PPCDSDCRDBUSIN[16], PPCDSDCRDBUSIN_OUT[16]);
buf B_PPCDSDCRDBUSIN17 (PPCDSDCRDBUSIN[17], PPCDSDCRDBUSIN_OUT[17]);
buf B_PPCDSDCRDBUSIN18 (PPCDSDCRDBUSIN[18], PPCDSDCRDBUSIN_OUT[18]);
buf B_PPCDSDCRDBUSIN19 (PPCDSDCRDBUSIN[19], PPCDSDCRDBUSIN_OUT[19]);
buf B_PPCDSDCRDBUSIN20 (PPCDSDCRDBUSIN[20], PPCDSDCRDBUSIN_OUT[20]);
buf B_PPCDSDCRDBUSIN21 (PPCDSDCRDBUSIN[21], PPCDSDCRDBUSIN_OUT[21]);
buf B_PPCDSDCRDBUSIN22 (PPCDSDCRDBUSIN[22], PPCDSDCRDBUSIN_OUT[22]);
buf B_PPCDSDCRDBUSIN23 (PPCDSDCRDBUSIN[23], PPCDSDCRDBUSIN_OUT[23]);
buf B_PPCDSDCRDBUSIN24 (PPCDSDCRDBUSIN[24], PPCDSDCRDBUSIN_OUT[24]);
buf B_PPCDSDCRDBUSIN25 (PPCDSDCRDBUSIN[25], PPCDSDCRDBUSIN_OUT[25]);
buf B_PPCDSDCRDBUSIN26 (PPCDSDCRDBUSIN[26], PPCDSDCRDBUSIN_OUT[26]);
buf B_PPCDSDCRDBUSIN27 (PPCDSDCRDBUSIN[27], PPCDSDCRDBUSIN_OUT[27]);
buf B_PPCDSDCRDBUSIN28 (PPCDSDCRDBUSIN[28], PPCDSDCRDBUSIN_OUT[28]);
buf B_PPCDSDCRDBUSIN29 (PPCDSDCRDBUSIN[29], PPCDSDCRDBUSIN_OUT[29]);
buf B_PPCDSDCRDBUSIN30 (PPCDSDCRDBUSIN[30], PPCDSDCRDBUSIN_OUT[30]);
buf B_PPCDSDCRDBUSIN31 (PPCDSDCRDBUSIN[31], PPCDSDCRDBUSIN_OUT[31]);
buf B_PPCEICINTERCONNECTIRQ (PPCEICINTERCONNECTIRQ, PPCEICINTERCONNECTIRQ_OUT);

buf B_PLBPPCS0RNW (PLBPPCS0RNW_IN, PLBPPCS0RNW);
buf B_PLBPPCS1RNW (PLBPPCS1RNW_IN, PLBPPCS1RNW);
buf B_CPMDCRCLK (CPMDCRCLK_IN, CPMDCRCLK);
buf B_CPMDMA0LLCLK (CPMDMA0LLCLK_IN, CPMDMA0LLCLK);
buf B_CPMDMA1LLCLK (CPMDMA1LLCLK_IN, CPMDMA1LLCLK);
buf B_CPMDMA2LLCLK (CPMDMA2LLCLK_IN, CPMDMA2LLCLK);
buf B_CPMDMA3LLCLK (CPMDMA3LLCLK_IN, CPMDMA3LLCLK);
buf B_CPMINTERCONNECTCLKNTO1 (CPMINTERCONNECTCLKNTO1_IN, CPMINTERCONNECTCLKNTO1);
buf B_CPMPPCMPLBCLK (CPMPPCMPLBCLK_IN, CPMPPCMPLBCLK);
buf B_CPMPPCS0PLBCLK (CPMPPCS0PLBCLK_IN, CPMPPCS0PLBCLK);
buf B_CPMPPCS1PLBCLK (CPMPPCS1PLBCLK_IN, CPMPPCS1PLBCLK);
buf B_DCRPPCDMACK (DCRPPCDMACK_IN, DCRPPCDMACK);
buf B_DCRPPCDMDBUSIN0 (DCRPPCDMDBUSIN_IN[0], DCRPPCDMDBUSIN[0]);
buf B_DCRPPCDMDBUSIN1 (DCRPPCDMDBUSIN_IN[1], DCRPPCDMDBUSIN[1]);
buf B_DCRPPCDMDBUSIN2 (DCRPPCDMDBUSIN_IN[2], DCRPPCDMDBUSIN[2]);
buf B_DCRPPCDMDBUSIN3 (DCRPPCDMDBUSIN_IN[3], DCRPPCDMDBUSIN[3]);
buf B_DCRPPCDMDBUSIN4 (DCRPPCDMDBUSIN_IN[4], DCRPPCDMDBUSIN[4]);
buf B_DCRPPCDMDBUSIN5 (DCRPPCDMDBUSIN_IN[5], DCRPPCDMDBUSIN[5]);
buf B_DCRPPCDMDBUSIN6 (DCRPPCDMDBUSIN_IN[6], DCRPPCDMDBUSIN[6]);
buf B_DCRPPCDMDBUSIN7 (DCRPPCDMDBUSIN_IN[7], DCRPPCDMDBUSIN[7]);
buf B_DCRPPCDMDBUSIN8 (DCRPPCDMDBUSIN_IN[8], DCRPPCDMDBUSIN[8]);
buf B_DCRPPCDMDBUSIN9 (DCRPPCDMDBUSIN_IN[9], DCRPPCDMDBUSIN[9]);
buf B_DCRPPCDMDBUSIN10 (DCRPPCDMDBUSIN_IN[10], DCRPPCDMDBUSIN[10]);
buf B_DCRPPCDMDBUSIN11 (DCRPPCDMDBUSIN_IN[11], DCRPPCDMDBUSIN[11]);
buf B_DCRPPCDMDBUSIN12 (DCRPPCDMDBUSIN_IN[12], DCRPPCDMDBUSIN[12]);
buf B_DCRPPCDMDBUSIN13 (DCRPPCDMDBUSIN_IN[13], DCRPPCDMDBUSIN[13]);
buf B_DCRPPCDMDBUSIN14 (DCRPPCDMDBUSIN_IN[14], DCRPPCDMDBUSIN[14]);
buf B_DCRPPCDMDBUSIN15 (DCRPPCDMDBUSIN_IN[15], DCRPPCDMDBUSIN[15]);
buf B_DCRPPCDMDBUSIN16 (DCRPPCDMDBUSIN_IN[16], DCRPPCDMDBUSIN[16]);
buf B_DCRPPCDMDBUSIN17 (DCRPPCDMDBUSIN_IN[17], DCRPPCDMDBUSIN[17]);
buf B_DCRPPCDMDBUSIN18 (DCRPPCDMDBUSIN_IN[18], DCRPPCDMDBUSIN[18]);
buf B_DCRPPCDMDBUSIN19 (DCRPPCDMDBUSIN_IN[19], DCRPPCDMDBUSIN[19]);
buf B_DCRPPCDMDBUSIN20 (DCRPPCDMDBUSIN_IN[20], DCRPPCDMDBUSIN[20]);
buf B_DCRPPCDMDBUSIN21 (DCRPPCDMDBUSIN_IN[21], DCRPPCDMDBUSIN[21]);
buf B_DCRPPCDMDBUSIN22 (DCRPPCDMDBUSIN_IN[22], DCRPPCDMDBUSIN[22]);
buf B_DCRPPCDMDBUSIN23 (DCRPPCDMDBUSIN_IN[23], DCRPPCDMDBUSIN[23]);
buf B_DCRPPCDMDBUSIN24 (DCRPPCDMDBUSIN_IN[24], DCRPPCDMDBUSIN[24]);
buf B_DCRPPCDMDBUSIN25 (DCRPPCDMDBUSIN_IN[25], DCRPPCDMDBUSIN[25]);
buf B_DCRPPCDMDBUSIN26 (DCRPPCDMDBUSIN_IN[26], DCRPPCDMDBUSIN[26]);
buf B_DCRPPCDMDBUSIN27 (DCRPPCDMDBUSIN_IN[27], DCRPPCDMDBUSIN[27]);
buf B_DCRPPCDMDBUSIN28 (DCRPPCDMDBUSIN_IN[28], DCRPPCDMDBUSIN[28]);
buf B_DCRPPCDMDBUSIN29 (DCRPPCDMDBUSIN_IN[29], DCRPPCDMDBUSIN[29]);
buf B_DCRPPCDMDBUSIN30 (DCRPPCDMDBUSIN_IN[30], DCRPPCDMDBUSIN[30]);
buf B_DCRPPCDMDBUSIN31 (DCRPPCDMDBUSIN_IN[31], DCRPPCDMDBUSIN[31]);
buf B_DCRPPCDMTIMEOUTWAIT (DCRPPCDMTIMEOUTWAIT_IN, DCRPPCDMTIMEOUTWAIT);
buf B_LLDMA0RSTENGINEREQ (LLDMA0RSTENGINEREQ_IN, LLDMA0RSTENGINEREQ);
buf B_LLDMA0RXD0 (LLDMA0RXD_IN[0], LLDMA0RXD[0]);
buf B_LLDMA0RXD1 (LLDMA0RXD_IN[1], LLDMA0RXD[1]);
buf B_LLDMA0RXD2 (LLDMA0RXD_IN[2], LLDMA0RXD[2]);
buf B_LLDMA0RXD3 (LLDMA0RXD_IN[3], LLDMA0RXD[3]);
buf B_LLDMA0RXD4 (LLDMA0RXD_IN[4], LLDMA0RXD[4]);
buf B_LLDMA0RXD5 (LLDMA0RXD_IN[5], LLDMA0RXD[5]);
buf B_LLDMA0RXD6 (LLDMA0RXD_IN[6], LLDMA0RXD[6]);
buf B_LLDMA0RXD7 (LLDMA0RXD_IN[7], LLDMA0RXD[7]);
buf B_LLDMA0RXD8 (LLDMA0RXD_IN[8], LLDMA0RXD[8]);
buf B_LLDMA0RXD9 (LLDMA0RXD_IN[9], LLDMA0RXD[9]);
buf B_LLDMA0RXD10 (LLDMA0RXD_IN[10], LLDMA0RXD[10]);
buf B_LLDMA0RXD11 (LLDMA0RXD_IN[11], LLDMA0RXD[11]);
buf B_LLDMA0RXD12 (LLDMA0RXD_IN[12], LLDMA0RXD[12]);
buf B_LLDMA0RXD13 (LLDMA0RXD_IN[13], LLDMA0RXD[13]);
buf B_LLDMA0RXD14 (LLDMA0RXD_IN[14], LLDMA0RXD[14]);
buf B_LLDMA0RXD15 (LLDMA0RXD_IN[15], LLDMA0RXD[15]);
buf B_LLDMA0RXD16 (LLDMA0RXD_IN[16], LLDMA0RXD[16]);
buf B_LLDMA0RXD17 (LLDMA0RXD_IN[17], LLDMA0RXD[17]);
buf B_LLDMA0RXD18 (LLDMA0RXD_IN[18], LLDMA0RXD[18]);
buf B_LLDMA0RXD19 (LLDMA0RXD_IN[19], LLDMA0RXD[19]);
buf B_LLDMA0RXD20 (LLDMA0RXD_IN[20], LLDMA0RXD[20]);
buf B_LLDMA0RXD21 (LLDMA0RXD_IN[21], LLDMA0RXD[21]);
buf B_LLDMA0RXD22 (LLDMA0RXD_IN[22], LLDMA0RXD[22]);
buf B_LLDMA0RXD23 (LLDMA0RXD_IN[23], LLDMA0RXD[23]);
buf B_LLDMA0RXD24 (LLDMA0RXD_IN[24], LLDMA0RXD[24]);
buf B_LLDMA0RXD25 (LLDMA0RXD_IN[25], LLDMA0RXD[25]);
buf B_LLDMA0RXD26 (LLDMA0RXD_IN[26], LLDMA0RXD[26]);
buf B_LLDMA0RXD27 (LLDMA0RXD_IN[27], LLDMA0RXD[27]);
buf B_LLDMA0RXD28 (LLDMA0RXD_IN[28], LLDMA0RXD[28]);
buf B_LLDMA0RXD29 (LLDMA0RXD_IN[29], LLDMA0RXD[29]);
buf B_LLDMA0RXD30 (LLDMA0RXD_IN[30], LLDMA0RXD[30]);
buf B_LLDMA0RXD31 (LLDMA0RXD_IN[31], LLDMA0RXD[31]);
buf B_LLDMA0RXEOFN (LLDMA0RXEOFN_IN, LLDMA0RXEOFN);
buf B_LLDMA0RXEOPN (LLDMA0RXEOPN_IN, LLDMA0RXEOPN);
buf B_LLDMA0RXREM0 (LLDMA0RXREM_IN[0], LLDMA0RXREM[0]);
buf B_LLDMA0RXREM1 (LLDMA0RXREM_IN[1], LLDMA0RXREM[1]);
buf B_LLDMA0RXREM2 (LLDMA0RXREM_IN[2], LLDMA0RXREM[2]);
buf B_LLDMA0RXREM3 (LLDMA0RXREM_IN[3], LLDMA0RXREM[3]);
buf B_LLDMA0RXSOFN (LLDMA0RXSOFN_IN, LLDMA0RXSOFN);
buf B_LLDMA0RXSOPN (LLDMA0RXSOPN_IN, LLDMA0RXSOPN);
buf B_LLDMA0RXSRCRDYN (LLDMA0RXSRCRDYN_IN, LLDMA0RXSRCRDYN);
buf B_LLDMA0TXDSTRDYN (LLDMA0TXDSTRDYN_IN, LLDMA0TXDSTRDYN);
buf B_LLDMA1RSTENGINEREQ (LLDMA1RSTENGINEREQ_IN, LLDMA1RSTENGINEREQ);
buf B_LLDMA1RXD0 (LLDMA1RXD_IN[0], LLDMA1RXD[0]);
buf B_LLDMA1RXD1 (LLDMA1RXD_IN[1], LLDMA1RXD[1]);
buf B_LLDMA1RXD2 (LLDMA1RXD_IN[2], LLDMA1RXD[2]);
buf B_LLDMA1RXD3 (LLDMA1RXD_IN[3], LLDMA1RXD[3]);
buf B_LLDMA1RXD4 (LLDMA1RXD_IN[4], LLDMA1RXD[4]);
buf B_LLDMA1RXD5 (LLDMA1RXD_IN[5], LLDMA1RXD[5]);
buf B_LLDMA1RXD6 (LLDMA1RXD_IN[6], LLDMA1RXD[6]);
buf B_LLDMA1RXD7 (LLDMA1RXD_IN[7], LLDMA1RXD[7]);
buf B_LLDMA1RXD8 (LLDMA1RXD_IN[8], LLDMA1RXD[8]);
buf B_LLDMA1RXD9 (LLDMA1RXD_IN[9], LLDMA1RXD[9]);
buf B_LLDMA1RXD10 (LLDMA1RXD_IN[10], LLDMA1RXD[10]);
buf B_LLDMA1RXD11 (LLDMA1RXD_IN[11], LLDMA1RXD[11]);
buf B_LLDMA1RXD12 (LLDMA1RXD_IN[12], LLDMA1RXD[12]);
buf B_LLDMA1RXD13 (LLDMA1RXD_IN[13], LLDMA1RXD[13]);
buf B_LLDMA1RXD14 (LLDMA1RXD_IN[14], LLDMA1RXD[14]);
buf B_LLDMA1RXD15 (LLDMA1RXD_IN[15], LLDMA1RXD[15]);
buf B_LLDMA1RXD16 (LLDMA1RXD_IN[16], LLDMA1RXD[16]);
buf B_LLDMA1RXD17 (LLDMA1RXD_IN[17], LLDMA1RXD[17]);
buf B_LLDMA1RXD18 (LLDMA1RXD_IN[18], LLDMA1RXD[18]);
buf B_LLDMA1RXD19 (LLDMA1RXD_IN[19], LLDMA1RXD[19]);
buf B_LLDMA1RXD20 (LLDMA1RXD_IN[20], LLDMA1RXD[20]);
buf B_LLDMA1RXD21 (LLDMA1RXD_IN[21], LLDMA1RXD[21]);
buf B_LLDMA1RXD22 (LLDMA1RXD_IN[22], LLDMA1RXD[22]);
buf B_LLDMA1RXD23 (LLDMA1RXD_IN[23], LLDMA1RXD[23]);
buf B_LLDMA1RXD24 (LLDMA1RXD_IN[24], LLDMA1RXD[24]);
buf B_LLDMA1RXD25 (LLDMA1RXD_IN[25], LLDMA1RXD[25]);
buf B_LLDMA1RXD26 (LLDMA1RXD_IN[26], LLDMA1RXD[26]);
buf B_LLDMA1RXD27 (LLDMA1RXD_IN[27], LLDMA1RXD[27]);
buf B_LLDMA1RXD28 (LLDMA1RXD_IN[28], LLDMA1RXD[28]);
buf B_LLDMA1RXD29 (LLDMA1RXD_IN[29], LLDMA1RXD[29]);
buf B_LLDMA1RXD30 (LLDMA1RXD_IN[30], LLDMA1RXD[30]);
buf B_LLDMA1RXD31 (LLDMA1RXD_IN[31], LLDMA1RXD[31]);
buf B_LLDMA1RXEOFN (LLDMA1RXEOFN_IN, LLDMA1RXEOFN);
buf B_LLDMA1RXEOPN (LLDMA1RXEOPN_IN, LLDMA1RXEOPN);
buf B_LLDMA1RXREM0 (LLDMA1RXREM_IN[0], LLDMA1RXREM[0]);
buf B_LLDMA1RXREM1 (LLDMA1RXREM_IN[1], LLDMA1RXREM[1]);
buf B_LLDMA1RXREM2 (LLDMA1RXREM_IN[2], LLDMA1RXREM[2]);
buf B_LLDMA1RXREM3 (LLDMA1RXREM_IN[3], LLDMA1RXREM[3]);
buf B_LLDMA1RXSOFN (LLDMA1RXSOFN_IN, LLDMA1RXSOFN);
buf B_LLDMA1RXSOPN (LLDMA1RXSOPN_IN, LLDMA1RXSOPN);
buf B_LLDMA1RXSRCRDYN (LLDMA1RXSRCRDYN_IN, LLDMA1RXSRCRDYN);
buf B_LLDMA1TXDSTRDYN (LLDMA1TXDSTRDYN_IN, LLDMA1TXDSTRDYN);
buf B_LLDMA2RSTENGINEREQ (LLDMA2RSTENGINEREQ_IN, LLDMA2RSTENGINEREQ);
buf B_LLDMA2RXD0 (LLDMA2RXD_IN[0], LLDMA2RXD[0]);
buf B_LLDMA2RXD1 (LLDMA2RXD_IN[1], LLDMA2RXD[1]);
buf B_LLDMA2RXD2 (LLDMA2RXD_IN[2], LLDMA2RXD[2]);
buf B_LLDMA2RXD3 (LLDMA2RXD_IN[3], LLDMA2RXD[3]);
buf B_LLDMA2RXD4 (LLDMA2RXD_IN[4], LLDMA2RXD[4]);
buf B_LLDMA2RXD5 (LLDMA2RXD_IN[5], LLDMA2RXD[5]);
buf B_LLDMA2RXD6 (LLDMA2RXD_IN[6], LLDMA2RXD[6]);
buf B_LLDMA2RXD7 (LLDMA2RXD_IN[7], LLDMA2RXD[7]);
buf B_LLDMA2RXD8 (LLDMA2RXD_IN[8], LLDMA2RXD[8]);
buf B_LLDMA2RXD9 (LLDMA2RXD_IN[9], LLDMA2RXD[9]);
buf B_LLDMA2RXD10 (LLDMA2RXD_IN[10], LLDMA2RXD[10]);
buf B_LLDMA2RXD11 (LLDMA2RXD_IN[11], LLDMA2RXD[11]);
buf B_LLDMA2RXD12 (LLDMA2RXD_IN[12], LLDMA2RXD[12]);
buf B_LLDMA2RXD13 (LLDMA2RXD_IN[13], LLDMA2RXD[13]);
buf B_LLDMA2RXD14 (LLDMA2RXD_IN[14], LLDMA2RXD[14]);
buf B_LLDMA2RXD15 (LLDMA2RXD_IN[15], LLDMA2RXD[15]);
buf B_LLDMA2RXD16 (LLDMA2RXD_IN[16], LLDMA2RXD[16]);
buf B_LLDMA2RXD17 (LLDMA2RXD_IN[17], LLDMA2RXD[17]);
buf B_LLDMA2RXD18 (LLDMA2RXD_IN[18], LLDMA2RXD[18]);
buf B_LLDMA2RXD19 (LLDMA2RXD_IN[19], LLDMA2RXD[19]);
buf B_LLDMA2RXD20 (LLDMA2RXD_IN[20], LLDMA2RXD[20]);
buf B_LLDMA2RXD21 (LLDMA2RXD_IN[21], LLDMA2RXD[21]);
buf B_LLDMA2RXD22 (LLDMA2RXD_IN[22], LLDMA2RXD[22]);
buf B_LLDMA2RXD23 (LLDMA2RXD_IN[23], LLDMA2RXD[23]);
buf B_LLDMA2RXD24 (LLDMA2RXD_IN[24], LLDMA2RXD[24]);
buf B_LLDMA2RXD25 (LLDMA2RXD_IN[25], LLDMA2RXD[25]);
buf B_LLDMA2RXD26 (LLDMA2RXD_IN[26], LLDMA2RXD[26]);
buf B_LLDMA2RXD27 (LLDMA2RXD_IN[27], LLDMA2RXD[27]);
buf B_LLDMA2RXD28 (LLDMA2RXD_IN[28], LLDMA2RXD[28]);
buf B_LLDMA2RXD29 (LLDMA2RXD_IN[29], LLDMA2RXD[29]);
buf B_LLDMA2RXD30 (LLDMA2RXD_IN[30], LLDMA2RXD[30]);
buf B_LLDMA2RXD31 (LLDMA2RXD_IN[31], LLDMA2RXD[31]);
buf B_LLDMA2RXEOFN (LLDMA2RXEOFN_IN, LLDMA2RXEOFN);
buf B_LLDMA2RXEOPN (LLDMA2RXEOPN_IN, LLDMA2RXEOPN);
buf B_LLDMA2RXREM0 (LLDMA2RXREM_IN[0], LLDMA2RXREM[0]);
buf B_LLDMA2RXREM1 (LLDMA2RXREM_IN[1], LLDMA2RXREM[1]);
buf B_LLDMA2RXREM2 (LLDMA2RXREM_IN[2], LLDMA2RXREM[2]);
buf B_LLDMA2RXREM3 (LLDMA2RXREM_IN[3], LLDMA2RXREM[3]);
buf B_LLDMA2RXSOFN (LLDMA2RXSOFN_IN, LLDMA2RXSOFN);
buf B_LLDMA2RXSOPN (LLDMA2RXSOPN_IN, LLDMA2RXSOPN);
buf B_LLDMA2RXSRCRDYN (LLDMA2RXSRCRDYN_IN, LLDMA2RXSRCRDYN);
buf B_LLDMA2TXDSTRDYN (LLDMA2TXDSTRDYN_IN, LLDMA2TXDSTRDYN);
buf B_LLDMA3RSTENGINEREQ (LLDMA3RSTENGINEREQ_IN, LLDMA3RSTENGINEREQ);
buf B_LLDMA3RXD0 (LLDMA3RXD_IN[0], LLDMA3RXD[0]);
buf B_LLDMA3RXD1 (LLDMA3RXD_IN[1], LLDMA3RXD[1]);
buf B_LLDMA3RXD2 (LLDMA3RXD_IN[2], LLDMA3RXD[2]);
buf B_LLDMA3RXD3 (LLDMA3RXD_IN[3], LLDMA3RXD[3]);
buf B_LLDMA3RXD4 (LLDMA3RXD_IN[4], LLDMA3RXD[4]);
buf B_LLDMA3RXD5 (LLDMA3RXD_IN[5], LLDMA3RXD[5]);
buf B_LLDMA3RXD6 (LLDMA3RXD_IN[6], LLDMA3RXD[6]);
buf B_LLDMA3RXD7 (LLDMA3RXD_IN[7], LLDMA3RXD[7]);
buf B_LLDMA3RXD8 (LLDMA3RXD_IN[8], LLDMA3RXD[8]);
buf B_LLDMA3RXD9 (LLDMA3RXD_IN[9], LLDMA3RXD[9]);
buf B_LLDMA3RXD10 (LLDMA3RXD_IN[10], LLDMA3RXD[10]);
buf B_LLDMA3RXD11 (LLDMA3RXD_IN[11], LLDMA3RXD[11]);
buf B_LLDMA3RXD12 (LLDMA3RXD_IN[12], LLDMA3RXD[12]);
buf B_LLDMA3RXD13 (LLDMA3RXD_IN[13], LLDMA3RXD[13]);
buf B_LLDMA3RXD14 (LLDMA3RXD_IN[14], LLDMA3RXD[14]);
buf B_LLDMA3RXD15 (LLDMA3RXD_IN[15], LLDMA3RXD[15]);
buf B_LLDMA3RXD16 (LLDMA3RXD_IN[16], LLDMA3RXD[16]);
buf B_LLDMA3RXD17 (LLDMA3RXD_IN[17], LLDMA3RXD[17]);
buf B_LLDMA3RXD18 (LLDMA3RXD_IN[18], LLDMA3RXD[18]);
buf B_LLDMA3RXD19 (LLDMA3RXD_IN[19], LLDMA3RXD[19]);
buf B_LLDMA3RXD20 (LLDMA3RXD_IN[20], LLDMA3RXD[20]);
buf B_LLDMA3RXD21 (LLDMA3RXD_IN[21], LLDMA3RXD[21]);
buf B_LLDMA3RXD22 (LLDMA3RXD_IN[22], LLDMA3RXD[22]);
buf B_LLDMA3RXD23 (LLDMA3RXD_IN[23], LLDMA3RXD[23]);
buf B_LLDMA3RXD24 (LLDMA3RXD_IN[24], LLDMA3RXD[24]);
buf B_LLDMA3RXD25 (LLDMA3RXD_IN[25], LLDMA3RXD[25]);
buf B_LLDMA3RXD26 (LLDMA3RXD_IN[26], LLDMA3RXD[26]);
buf B_LLDMA3RXD27 (LLDMA3RXD_IN[27], LLDMA3RXD[27]);
buf B_LLDMA3RXD28 (LLDMA3RXD_IN[28], LLDMA3RXD[28]);
buf B_LLDMA3RXD29 (LLDMA3RXD_IN[29], LLDMA3RXD[29]);
buf B_LLDMA3RXD30 (LLDMA3RXD_IN[30], LLDMA3RXD[30]);
buf B_LLDMA3RXD31 (LLDMA3RXD_IN[31], LLDMA3RXD[31]);
buf B_LLDMA3RXEOFN (LLDMA3RXEOFN_IN, LLDMA3RXEOFN);
buf B_LLDMA3RXEOPN (LLDMA3RXEOPN_IN, LLDMA3RXEOPN);
buf B_LLDMA3RXREM0 (LLDMA3RXREM_IN[0], LLDMA3RXREM[0]);
buf B_LLDMA3RXREM1 (LLDMA3RXREM_IN[1], LLDMA3RXREM[1]);
buf B_LLDMA3RXREM2 (LLDMA3RXREM_IN[2], LLDMA3RXREM[2]);
buf B_LLDMA3RXREM3 (LLDMA3RXREM_IN[3], LLDMA3RXREM[3]);
buf B_LLDMA3RXSOFN (LLDMA3RXSOFN_IN, LLDMA3RXSOFN);
buf B_LLDMA3RXSOPN (LLDMA3RXSOPN_IN, LLDMA3RXSOPN);
buf B_LLDMA3RXSRCRDYN (LLDMA3RXSRCRDYN_IN, LLDMA3RXSRCRDYN);
buf B_LLDMA3TXDSTRDYN (LLDMA3TXDSTRDYN_IN, LLDMA3TXDSTRDYN);
buf B_PLBPPCMADDRACK (PLBPPCMADDRACK_IN, PLBPPCMADDRACK);
buf B_PLBPPCMMBUSY (PLBPPCMMBUSY_IN, PLBPPCMMBUSY);
buf B_PLBPPCMMIRQ (PLBPPCMMIRQ_IN, PLBPPCMMIRQ);
buf B_PLBPPCMMRDERR (PLBPPCMMRDERR_IN, PLBPPCMMRDERR);
buf B_PLBPPCMMWRERR (PLBPPCMMWRERR_IN, PLBPPCMMWRERR);
buf B_PLBPPCMRDBTERM (PLBPPCMRDBTERM_IN, PLBPPCMRDBTERM);
buf B_PLBPPCMRDDACK (PLBPPCMRDDACK_IN, PLBPPCMRDDACK);
buf B_PLBPPCMRDDBUS0 (PLBPPCMRDDBUS_IN[0], PLBPPCMRDDBUS[0]);
buf B_PLBPPCMRDDBUS1 (PLBPPCMRDDBUS_IN[1], PLBPPCMRDDBUS[1]);
buf B_PLBPPCMRDDBUS2 (PLBPPCMRDDBUS_IN[2], PLBPPCMRDDBUS[2]);
buf B_PLBPPCMRDDBUS3 (PLBPPCMRDDBUS_IN[3], PLBPPCMRDDBUS[3]);
buf B_PLBPPCMRDDBUS4 (PLBPPCMRDDBUS_IN[4], PLBPPCMRDDBUS[4]);
buf B_PLBPPCMRDDBUS5 (PLBPPCMRDDBUS_IN[5], PLBPPCMRDDBUS[5]);
buf B_PLBPPCMRDDBUS6 (PLBPPCMRDDBUS_IN[6], PLBPPCMRDDBUS[6]);
buf B_PLBPPCMRDDBUS7 (PLBPPCMRDDBUS_IN[7], PLBPPCMRDDBUS[7]);
buf B_PLBPPCMRDDBUS8 (PLBPPCMRDDBUS_IN[8], PLBPPCMRDDBUS[8]);
buf B_PLBPPCMRDDBUS9 (PLBPPCMRDDBUS_IN[9], PLBPPCMRDDBUS[9]);
buf B_PLBPPCMRDDBUS10 (PLBPPCMRDDBUS_IN[10], PLBPPCMRDDBUS[10]);
buf B_PLBPPCMRDDBUS11 (PLBPPCMRDDBUS_IN[11], PLBPPCMRDDBUS[11]);
buf B_PLBPPCMRDDBUS12 (PLBPPCMRDDBUS_IN[12], PLBPPCMRDDBUS[12]);
buf B_PLBPPCMRDDBUS13 (PLBPPCMRDDBUS_IN[13], PLBPPCMRDDBUS[13]);
buf B_PLBPPCMRDDBUS14 (PLBPPCMRDDBUS_IN[14], PLBPPCMRDDBUS[14]);
buf B_PLBPPCMRDDBUS15 (PLBPPCMRDDBUS_IN[15], PLBPPCMRDDBUS[15]);
buf B_PLBPPCMRDDBUS16 (PLBPPCMRDDBUS_IN[16], PLBPPCMRDDBUS[16]);
buf B_PLBPPCMRDDBUS17 (PLBPPCMRDDBUS_IN[17], PLBPPCMRDDBUS[17]);
buf B_PLBPPCMRDDBUS18 (PLBPPCMRDDBUS_IN[18], PLBPPCMRDDBUS[18]);
buf B_PLBPPCMRDDBUS19 (PLBPPCMRDDBUS_IN[19], PLBPPCMRDDBUS[19]);
buf B_PLBPPCMRDDBUS20 (PLBPPCMRDDBUS_IN[20], PLBPPCMRDDBUS[20]);
buf B_PLBPPCMRDDBUS21 (PLBPPCMRDDBUS_IN[21], PLBPPCMRDDBUS[21]);
buf B_PLBPPCMRDDBUS22 (PLBPPCMRDDBUS_IN[22], PLBPPCMRDDBUS[22]);
buf B_PLBPPCMRDDBUS23 (PLBPPCMRDDBUS_IN[23], PLBPPCMRDDBUS[23]);
buf B_PLBPPCMRDDBUS24 (PLBPPCMRDDBUS_IN[24], PLBPPCMRDDBUS[24]);
buf B_PLBPPCMRDDBUS25 (PLBPPCMRDDBUS_IN[25], PLBPPCMRDDBUS[25]);
buf B_PLBPPCMRDDBUS26 (PLBPPCMRDDBUS_IN[26], PLBPPCMRDDBUS[26]);
buf B_PLBPPCMRDDBUS27 (PLBPPCMRDDBUS_IN[27], PLBPPCMRDDBUS[27]);
buf B_PLBPPCMRDDBUS28 (PLBPPCMRDDBUS_IN[28], PLBPPCMRDDBUS[28]);
buf B_PLBPPCMRDDBUS29 (PLBPPCMRDDBUS_IN[29], PLBPPCMRDDBUS[29]);
buf B_PLBPPCMRDDBUS30 (PLBPPCMRDDBUS_IN[30], PLBPPCMRDDBUS[30]);
buf B_PLBPPCMRDDBUS31 (PLBPPCMRDDBUS_IN[31], PLBPPCMRDDBUS[31]);
buf B_PLBPPCMRDDBUS32 (PLBPPCMRDDBUS_IN[32], PLBPPCMRDDBUS[32]);
buf B_PLBPPCMRDDBUS33 (PLBPPCMRDDBUS_IN[33], PLBPPCMRDDBUS[33]);
buf B_PLBPPCMRDDBUS34 (PLBPPCMRDDBUS_IN[34], PLBPPCMRDDBUS[34]);
buf B_PLBPPCMRDDBUS35 (PLBPPCMRDDBUS_IN[35], PLBPPCMRDDBUS[35]);
buf B_PLBPPCMRDDBUS36 (PLBPPCMRDDBUS_IN[36], PLBPPCMRDDBUS[36]);
buf B_PLBPPCMRDDBUS37 (PLBPPCMRDDBUS_IN[37], PLBPPCMRDDBUS[37]);
buf B_PLBPPCMRDDBUS38 (PLBPPCMRDDBUS_IN[38], PLBPPCMRDDBUS[38]);
buf B_PLBPPCMRDDBUS39 (PLBPPCMRDDBUS_IN[39], PLBPPCMRDDBUS[39]);
buf B_PLBPPCMRDDBUS40 (PLBPPCMRDDBUS_IN[40], PLBPPCMRDDBUS[40]);
buf B_PLBPPCMRDDBUS41 (PLBPPCMRDDBUS_IN[41], PLBPPCMRDDBUS[41]);
buf B_PLBPPCMRDDBUS42 (PLBPPCMRDDBUS_IN[42], PLBPPCMRDDBUS[42]);
buf B_PLBPPCMRDDBUS43 (PLBPPCMRDDBUS_IN[43], PLBPPCMRDDBUS[43]);
buf B_PLBPPCMRDDBUS44 (PLBPPCMRDDBUS_IN[44], PLBPPCMRDDBUS[44]);
buf B_PLBPPCMRDDBUS45 (PLBPPCMRDDBUS_IN[45], PLBPPCMRDDBUS[45]);
buf B_PLBPPCMRDDBUS46 (PLBPPCMRDDBUS_IN[46], PLBPPCMRDDBUS[46]);
buf B_PLBPPCMRDDBUS47 (PLBPPCMRDDBUS_IN[47], PLBPPCMRDDBUS[47]);
buf B_PLBPPCMRDDBUS48 (PLBPPCMRDDBUS_IN[48], PLBPPCMRDDBUS[48]);
buf B_PLBPPCMRDDBUS49 (PLBPPCMRDDBUS_IN[49], PLBPPCMRDDBUS[49]);
buf B_PLBPPCMRDDBUS50 (PLBPPCMRDDBUS_IN[50], PLBPPCMRDDBUS[50]);
buf B_PLBPPCMRDDBUS51 (PLBPPCMRDDBUS_IN[51], PLBPPCMRDDBUS[51]);
buf B_PLBPPCMRDDBUS52 (PLBPPCMRDDBUS_IN[52], PLBPPCMRDDBUS[52]);
buf B_PLBPPCMRDDBUS53 (PLBPPCMRDDBUS_IN[53], PLBPPCMRDDBUS[53]);
buf B_PLBPPCMRDDBUS54 (PLBPPCMRDDBUS_IN[54], PLBPPCMRDDBUS[54]);
buf B_PLBPPCMRDDBUS55 (PLBPPCMRDDBUS_IN[55], PLBPPCMRDDBUS[55]);
buf B_PLBPPCMRDDBUS56 (PLBPPCMRDDBUS_IN[56], PLBPPCMRDDBUS[56]);
buf B_PLBPPCMRDDBUS57 (PLBPPCMRDDBUS_IN[57], PLBPPCMRDDBUS[57]);
buf B_PLBPPCMRDDBUS58 (PLBPPCMRDDBUS_IN[58], PLBPPCMRDDBUS[58]);
buf B_PLBPPCMRDDBUS59 (PLBPPCMRDDBUS_IN[59], PLBPPCMRDDBUS[59]);
buf B_PLBPPCMRDDBUS60 (PLBPPCMRDDBUS_IN[60], PLBPPCMRDDBUS[60]);
buf B_PLBPPCMRDDBUS61 (PLBPPCMRDDBUS_IN[61], PLBPPCMRDDBUS[61]);
buf B_PLBPPCMRDDBUS62 (PLBPPCMRDDBUS_IN[62], PLBPPCMRDDBUS[62]);
buf B_PLBPPCMRDDBUS63 (PLBPPCMRDDBUS_IN[63], PLBPPCMRDDBUS[63]);
buf B_PLBPPCMRDDBUS64 (PLBPPCMRDDBUS_IN[64], PLBPPCMRDDBUS[64]);
buf B_PLBPPCMRDDBUS65 (PLBPPCMRDDBUS_IN[65], PLBPPCMRDDBUS[65]);
buf B_PLBPPCMRDDBUS66 (PLBPPCMRDDBUS_IN[66], PLBPPCMRDDBUS[66]);
buf B_PLBPPCMRDDBUS67 (PLBPPCMRDDBUS_IN[67], PLBPPCMRDDBUS[67]);
buf B_PLBPPCMRDDBUS68 (PLBPPCMRDDBUS_IN[68], PLBPPCMRDDBUS[68]);
buf B_PLBPPCMRDDBUS69 (PLBPPCMRDDBUS_IN[69], PLBPPCMRDDBUS[69]);
buf B_PLBPPCMRDDBUS70 (PLBPPCMRDDBUS_IN[70], PLBPPCMRDDBUS[70]);
buf B_PLBPPCMRDDBUS71 (PLBPPCMRDDBUS_IN[71], PLBPPCMRDDBUS[71]);
buf B_PLBPPCMRDDBUS72 (PLBPPCMRDDBUS_IN[72], PLBPPCMRDDBUS[72]);
buf B_PLBPPCMRDDBUS73 (PLBPPCMRDDBUS_IN[73], PLBPPCMRDDBUS[73]);
buf B_PLBPPCMRDDBUS74 (PLBPPCMRDDBUS_IN[74], PLBPPCMRDDBUS[74]);
buf B_PLBPPCMRDDBUS75 (PLBPPCMRDDBUS_IN[75], PLBPPCMRDDBUS[75]);
buf B_PLBPPCMRDDBUS76 (PLBPPCMRDDBUS_IN[76], PLBPPCMRDDBUS[76]);
buf B_PLBPPCMRDDBUS77 (PLBPPCMRDDBUS_IN[77], PLBPPCMRDDBUS[77]);
buf B_PLBPPCMRDDBUS78 (PLBPPCMRDDBUS_IN[78], PLBPPCMRDDBUS[78]);
buf B_PLBPPCMRDDBUS79 (PLBPPCMRDDBUS_IN[79], PLBPPCMRDDBUS[79]);
buf B_PLBPPCMRDDBUS80 (PLBPPCMRDDBUS_IN[80], PLBPPCMRDDBUS[80]);
buf B_PLBPPCMRDDBUS81 (PLBPPCMRDDBUS_IN[81], PLBPPCMRDDBUS[81]);
buf B_PLBPPCMRDDBUS82 (PLBPPCMRDDBUS_IN[82], PLBPPCMRDDBUS[82]);
buf B_PLBPPCMRDDBUS83 (PLBPPCMRDDBUS_IN[83], PLBPPCMRDDBUS[83]);
buf B_PLBPPCMRDDBUS84 (PLBPPCMRDDBUS_IN[84], PLBPPCMRDDBUS[84]);
buf B_PLBPPCMRDDBUS85 (PLBPPCMRDDBUS_IN[85], PLBPPCMRDDBUS[85]);
buf B_PLBPPCMRDDBUS86 (PLBPPCMRDDBUS_IN[86], PLBPPCMRDDBUS[86]);
buf B_PLBPPCMRDDBUS87 (PLBPPCMRDDBUS_IN[87], PLBPPCMRDDBUS[87]);
buf B_PLBPPCMRDDBUS88 (PLBPPCMRDDBUS_IN[88], PLBPPCMRDDBUS[88]);
buf B_PLBPPCMRDDBUS89 (PLBPPCMRDDBUS_IN[89], PLBPPCMRDDBUS[89]);
buf B_PLBPPCMRDDBUS90 (PLBPPCMRDDBUS_IN[90], PLBPPCMRDDBUS[90]);
buf B_PLBPPCMRDDBUS91 (PLBPPCMRDDBUS_IN[91], PLBPPCMRDDBUS[91]);
buf B_PLBPPCMRDDBUS92 (PLBPPCMRDDBUS_IN[92], PLBPPCMRDDBUS[92]);
buf B_PLBPPCMRDDBUS93 (PLBPPCMRDDBUS_IN[93], PLBPPCMRDDBUS[93]);
buf B_PLBPPCMRDDBUS94 (PLBPPCMRDDBUS_IN[94], PLBPPCMRDDBUS[94]);
buf B_PLBPPCMRDDBUS95 (PLBPPCMRDDBUS_IN[95], PLBPPCMRDDBUS[95]);
buf B_PLBPPCMRDDBUS96 (PLBPPCMRDDBUS_IN[96], PLBPPCMRDDBUS[96]);
buf B_PLBPPCMRDDBUS97 (PLBPPCMRDDBUS_IN[97], PLBPPCMRDDBUS[97]);
buf B_PLBPPCMRDDBUS98 (PLBPPCMRDDBUS_IN[98], PLBPPCMRDDBUS[98]);
buf B_PLBPPCMRDDBUS99 (PLBPPCMRDDBUS_IN[99], PLBPPCMRDDBUS[99]);
buf B_PLBPPCMRDDBUS100 (PLBPPCMRDDBUS_IN[100], PLBPPCMRDDBUS[100]);
buf B_PLBPPCMRDDBUS101 (PLBPPCMRDDBUS_IN[101], PLBPPCMRDDBUS[101]);
buf B_PLBPPCMRDDBUS102 (PLBPPCMRDDBUS_IN[102], PLBPPCMRDDBUS[102]);
buf B_PLBPPCMRDDBUS103 (PLBPPCMRDDBUS_IN[103], PLBPPCMRDDBUS[103]);
buf B_PLBPPCMRDDBUS104 (PLBPPCMRDDBUS_IN[104], PLBPPCMRDDBUS[104]);
buf B_PLBPPCMRDDBUS105 (PLBPPCMRDDBUS_IN[105], PLBPPCMRDDBUS[105]);
buf B_PLBPPCMRDDBUS106 (PLBPPCMRDDBUS_IN[106], PLBPPCMRDDBUS[106]);
buf B_PLBPPCMRDDBUS107 (PLBPPCMRDDBUS_IN[107], PLBPPCMRDDBUS[107]);
buf B_PLBPPCMRDDBUS108 (PLBPPCMRDDBUS_IN[108], PLBPPCMRDDBUS[108]);
buf B_PLBPPCMRDDBUS109 (PLBPPCMRDDBUS_IN[109], PLBPPCMRDDBUS[109]);
buf B_PLBPPCMRDDBUS110 (PLBPPCMRDDBUS_IN[110], PLBPPCMRDDBUS[110]);
buf B_PLBPPCMRDDBUS111 (PLBPPCMRDDBUS_IN[111], PLBPPCMRDDBUS[111]);
buf B_PLBPPCMRDDBUS112 (PLBPPCMRDDBUS_IN[112], PLBPPCMRDDBUS[112]);
buf B_PLBPPCMRDDBUS113 (PLBPPCMRDDBUS_IN[113], PLBPPCMRDDBUS[113]);
buf B_PLBPPCMRDDBUS114 (PLBPPCMRDDBUS_IN[114], PLBPPCMRDDBUS[114]);
buf B_PLBPPCMRDDBUS115 (PLBPPCMRDDBUS_IN[115], PLBPPCMRDDBUS[115]);
buf B_PLBPPCMRDDBUS116 (PLBPPCMRDDBUS_IN[116], PLBPPCMRDDBUS[116]);
buf B_PLBPPCMRDDBUS117 (PLBPPCMRDDBUS_IN[117], PLBPPCMRDDBUS[117]);
buf B_PLBPPCMRDDBUS118 (PLBPPCMRDDBUS_IN[118], PLBPPCMRDDBUS[118]);
buf B_PLBPPCMRDDBUS119 (PLBPPCMRDDBUS_IN[119], PLBPPCMRDDBUS[119]);
buf B_PLBPPCMRDDBUS120 (PLBPPCMRDDBUS_IN[120], PLBPPCMRDDBUS[120]);
buf B_PLBPPCMRDDBUS121 (PLBPPCMRDDBUS_IN[121], PLBPPCMRDDBUS[121]);
buf B_PLBPPCMRDDBUS122 (PLBPPCMRDDBUS_IN[122], PLBPPCMRDDBUS[122]);
buf B_PLBPPCMRDDBUS123 (PLBPPCMRDDBUS_IN[123], PLBPPCMRDDBUS[123]);
buf B_PLBPPCMRDDBUS124 (PLBPPCMRDDBUS_IN[124], PLBPPCMRDDBUS[124]);
buf B_PLBPPCMRDDBUS125 (PLBPPCMRDDBUS_IN[125], PLBPPCMRDDBUS[125]);
buf B_PLBPPCMRDDBUS126 (PLBPPCMRDDBUS_IN[126], PLBPPCMRDDBUS[126]);
buf B_PLBPPCMRDDBUS127 (PLBPPCMRDDBUS_IN[127], PLBPPCMRDDBUS[127]);
buf B_PLBPPCMRDPENDPRI0 (PLBPPCMRDPENDPRI_IN[0], PLBPPCMRDPENDPRI[0]);
buf B_PLBPPCMRDPENDPRI1 (PLBPPCMRDPENDPRI_IN[1], PLBPPCMRDPENDPRI[1]);
buf B_PLBPPCMRDPENDREQ (PLBPPCMRDPENDREQ_IN, PLBPPCMRDPENDREQ);
buf B_PLBPPCMRDWDADDR0 (PLBPPCMRDWDADDR_IN[0], PLBPPCMRDWDADDR[0]);
buf B_PLBPPCMRDWDADDR1 (PLBPPCMRDWDADDR_IN[1], PLBPPCMRDWDADDR[1]);
buf B_PLBPPCMRDWDADDR2 (PLBPPCMRDWDADDR_IN[2], PLBPPCMRDWDADDR[2]);
buf B_PLBPPCMRDWDADDR3 (PLBPPCMRDWDADDR_IN[3], PLBPPCMRDWDADDR[3]);
buf B_PLBPPCMREARBITRATE (PLBPPCMREARBITRATE_IN, PLBPPCMREARBITRATE);
buf B_PLBPPCMREQPRI0 (PLBPPCMREQPRI_IN[0], PLBPPCMREQPRI[0]);
buf B_PLBPPCMREQPRI1 (PLBPPCMREQPRI_IN[1], PLBPPCMREQPRI[1]);
buf B_PLBPPCMSSIZE0 (PLBPPCMSSIZE_IN[0], PLBPPCMSSIZE[0]);
buf B_PLBPPCMSSIZE1 (PLBPPCMSSIZE_IN[1], PLBPPCMSSIZE[1]);
buf B_PLBPPCMTIMEOUT (PLBPPCMTIMEOUT_IN, PLBPPCMTIMEOUT);
buf B_PLBPPCMWRBTERM (PLBPPCMWRBTERM_IN, PLBPPCMWRBTERM);
buf B_PLBPPCMWRDACK (PLBPPCMWRDACK_IN, PLBPPCMWRDACK);
buf B_PLBPPCMWRPENDPRI0 (PLBPPCMWRPENDPRI_IN[0], PLBPPCMWRPENDPRI[0]);
buf B_PLBPPCMWRPENDPRI1 (PLBPPCMWRPENDPRI_IN[1], PLBPPCMWRPENDPRI[1]);
buf B_PLBPPCMWRPENDREQ (PLBPPCMWRPENDREQ_IN, PLBPPCMWRPENDREQ);
buf B_PLBPPCS0ABORT (PLBPPCS0ABORT_IN, PLBPPCS0ABORT);
buf B_PLBPPCS0ABUS0 (PLBPPCS0ABUS_IN[0], PLBPPCS0ABUS[0]);
buf B_PLBPPCS0ABUS1 (PLBPPCS0ABUS_IN[1], PLBPPCS0ABUS[1]);
buf B_PLBPPCS0ABUS2 (PLBPPCS0ABUS_IN[2], PLBPPCS0ABUS[2]);
buf B_PLBPPCS0ABUS3 (PLBPPCS0ABUS_IN[3], PLBPPCS0ABUS[3]);
buf B_PLBPPCS0ABUS4 (PLBPPCS0ABUS_IN[4], PLBPPCS0ABUS[4]);
buf B_PLBPPCS0ABUS5 (PLBPPCS0ABUS_IN[5], PLBPPCS0ABUS[5]);
buf B_PLBPPCS0ABUS6 (PLBPPCS0ABUS_IN[6], PLBPPCS0ABUS[6]);
buf B_PLBPPCS0ABUS7 (PLBPPCS0ABUS_IN[7], PLBPPCS0ABUS[7]);
buf B_PLBPPCS0ABUS8 (PLBPPCS0ABUS_IN[8], PLBPPCS0ABUS[8]);
buf B_PLBPPCS0ABUS9 (PLBPPCS0ABUS_IN[9], PLBPPCS0ABUS[9]);
buf B_PLBPPCS0ABUS10 (PLBPPCS0ABUS_IN[10], PLBPPCS0ABUS[10]);
buf B_PLBPPCS0ABUS11 (PLBPPCS0ABUS_IN[11], PLBPPCS0ABUS[11]);
buf B_PLBPPCS0ABUS12 (PLBPPCS0ABUS_IN[12], PLBPPCS0ABUS[12]);
buf B_PLBPPCS0ABUS13 (PLBPPCS0ABUS_IN[13], PLBPPCS0ABUS[13]);
buf B_PLBPPCS0ABUS14 (PLBPPCS0ABUS_IN[14], PLBPPCS0ABUS[14]);
buf B_PLBPPCS0ABUS15 (PLBPPCS0ABUS_IN[15], PLBPPCS0ABUS[15]);
buf B_PLBPPCS0ABUS16 (PLBPPCS0ABUS_IN[16], PLBPPCS0ABUS[16]);
buf B_PLBPPCS0ABUS17 (PLBPPCS0ABUS_IN[17], PLBPPCS0ABUS[17]);
buf B_PLBPPCS0ABUS18 (PLBPPCS0ABUS_IN[18], PLBPPCS0ABUS[18]);
buf B_PLBPPCS0ABUS19 (PLBPPCS0ABUS_IN[19], PLBPPCS0ABUS[19]);
buf B_PLBPPCS0ABUS20 (PLBPPCS0ABUS_IN[20], PLBPPCS0ABUS[20]);
buf B_PLBPPCS0ABUS21 (PLBPPCS0ABUS_IN[21], PLBPPCS0ABUS[21]);
buf B_PLBPPCS0ABUS22 (PLBPPCS0ABUS_IN[22], PLBPPCS0ABUS[22]);
buf B_PLBPPCS0ABUS23 (PLBPPCS0ABUS_IN[23], PLBPPCS0ABUS[23]);
buf B_PLBPPCS0ABUS24 (PLBPPCS0ABUS_IN[24], PLBPPCS0ABUS[24]);
buf B_PLBPPCS0ABUS25 (PLBPPCS0ABUS_IN[25], PLBPPCS0ABUS[25]);
buf B_PLBPPCS0ABUS26 (PLBPPCS0ABUS_IN[26], PLBPPCS0ABUS[26]);
buf B_PLBPPCS0ABUS27 (PLBPPCS0ABUS_IN[27], PLBPPCS0ABUS[27]);
buf B_PLBPPCS0ABUS28 (PLBPPCS0ABUS_IN[28], PLBPPCS0ABUS[28]);
buf B_PLBPPCS0ABUS29 (PLBPPCS0ABUS_IN[29], PLBPPCS0ABUS[29]);
buf B_PLBPPCS0ABUS30 (PLBPPCS0ABUS_IN[30], PLBPPCS0ABUS[30]);
buf B_PLBPPCS0ABUS31 (PLBPPCS0ABUS_IN[31], PLBPPCS0ABUS[31]);
buf B_PLBPPCS0BE0 (PLBPPCS0BE_IN[0], PLBPPCS0BE[0]);
buf B_PLBPPCS0BE1 (PLBPPCS0BE_IN[1], PLBPPCS0BE[1]);
buf B_PLBPPCS0BE2 (PLBPPCS0BE_IN[2], PLBPPCS0BE[2]);
buf B_PLBPPCS0BE3 (PLBPPCS0BE_IN[3], PLBPPCS0BE[3]);
buf B_PLBPPCS0BE4 (PLBPPCS0BE_IN[4], PLBPPCS0BE[4]);
buf B_PLBPPCS0BE5 (PLBPPCS0BE_IN[5], PLBPPCS0BE[5]);
buf B_PLBPPCS0BE6 (PLBPPCS0BE_IN[6], PLBPPCS0BE[6]);
buf B_PLBPPCS0BE7 (PLBPPCS0BE_IN[7], PLBPPCS0BE[7]);
buf B_PLBPPCS0BE8 (PLBPPCS0BE_IN[8], PLBPPCS0BE[8]);
buf B_PLBPPCS0BE9 (PLBPPCS0BE_IN[9], PLBPPCS0BE[9]);
buf B_PLBPPCS0BE10 (PLBPPCS0BE_IN[10], PLBPPCS0BE[10]);
buf B_PLBPPCS0BE11 (PLBPPCS0BE_IN[11], PLBPPCS0BE[11]);
buf B_PLBPPCS0BE12 (PLBPPCS0BE_IN[12], PLBPPCS0BE[12]);
buf B_PLBPPCS0BE13 (PLBPPCS0BE_IN[13], PLBPPCS0BE[13]);
buf B_PLBPPCS0BE14 (PLBPPCS0BE_IN[14], PLBPPCS0BE[14]);
buf B_PLBPPCS0BE15 (PLBPPCS0BE_IN[15], PLBPPCS0BE[15]);
buf B_PLBPPCS0BUSLOCK (PLBPPCS0BUSLOCK_IN, PLBPPCS0BUSLOCK);
buf B_PLBPPCS0LOCKERR (PLBPPCS0LOCKERR_IN, PLBPPCS0LOCKERR);
buf B_PLBPPCS0MASTERID0 (PLBPPCS0MASTERID_IN[0], PLBPPCS0MASTERID[0]);
buf B_PLBPPCS0MASTERID1 (PLBPPCS0MASTERID_IN[1], PLBPPCS0MASTERID[1]);
buf B_PLBPPCS0MSIZE0 (PLBPPCS0MSIZE_IN[0], PLBPPCS0MSIZE[0]);
buf B_PLBPPCS0MSIZE1 (PLBPPCS0MSIZE_IN[1], PLBPPCS0MSIZE[1]);
buf B_PLBPPCS0PAVALID (PLBPPCS0PAVALID_IN, PLBPPCS0PAVALID);
buf B_PLBPPCS0RDBURST (PLBPPCS0RDBURST_IN, PLBPPCS0RDBURST);
buf B_PLBPPCS0RDPENDPRI0 (PLBPPCS0RDPENDPRI_IN[0], PLBPPCS0RDPENDPRI[0]);
buf B_PLBPPCS0RDPENDPRI1 (PLBPPCS0RDPENDPRI_IN[1], PLBPPCS0RDPENDPRI[1]);
buf B_PLBPPCS0RDPENDREQ (PLBPPCS0RDPENDREQ_IN, PLBPPCS0RDPENDREQ);
buf B_PLBPPCS0RDPRIM (PLBPPCS0RDPRIM_IN, PLBPPCS0RDPRIM);
buf B_PLBPPCS0REQPRI0 (PLBPPCS0REQPRI_IN[0], PLBPPCS0REQPRI[0]);
buf B_PLBPPCS0REQPRI1 (PLBPPCS0REQPRI_IN[1], PLBPPCS0REQPRI[1]);
buf B_PLBPPCS0SAVALID (PLBPPCS0SAVALID_IN, PLBPPCS0SAVALID);
buf B_PLBPPCS0SIZE0 (PLBPPCS0SIZE_IN[0], PLBPPCS0SIZE[0]);
buf B_PLBPPCS0SIZE1 (PLBPPCS0SIZE_IN[1], PLBPPCS0SIZE[1]);
buf B_PLBPPCS0SIZE2 (PLBPPCS0SIZE_IN[2], PLBPPCS0SIZE[2]);
buf B_PLBPPCS0SIZE3 (PLBPPCS0SIZE_IN[3], PLBPPCS0SIZE[3]);
buf B_PLBPPCS0TATTRIBUTE0 (PLBPPCS0TATTRIBUTE_IN[0], PLBPPCS0TATTRIBUTE[0]);
buf B_PLBPPCS0TATTRIBUTE1 (PLBPPCS0TATTRIBUTE_IN[1], PLBPPCS0TATTRIBUTE[1]);
buf B_PLBPPCS0TATTRIBUTE2 (PLBPPCS0TATTRIBUTE_IN[2], PLBPPCS0TATTRIBUTE[2]);
buf B_PLBPPCS0TATTRIBUTE3 (PLBPPCS0TATTRIBUTE_IN[3], PLBPPCS0TATTRIBUTE[3]);
buf B_PLBPPCS0TATTRIBUTE4 (PLBPPCS0TATTRIBUTE_IN[4], PLBPPCS0TATTRIBUTE[4]);
buf B_PLBPPCS0TATTRIBUTE5 (PLBPPCS0TATTRIBUTE_IN[5], PLBPPCS0TATTRIBUTE[5]);
buf B_PLBPPCS0TATTRIBUTE6 (PLBPPCS0TATTRIBUTE_IN[6], PLBPPCS0TATTRIBUTE[6]);
buf B_PLBPPCS0TATTRIBUTE7 (PLBPPCS0TATTRIBUTE_IN[7], PLBPPCS0TATTRIBUTE[7]);
buf B_PLBPPCS0TATTRIBUTE8 (PLBPPCS0TATTRIBUTE_IN[8], PLBPPCS0TATTRIBUTE[8]);
buf B_PLBPPCS0TATTRIBUTE9 (PLBPPCS0TATTRIBUTE_IN[9], PLBPPCS0TATTRIBUTE[9]);
buf B_PLBPPCS0TATTRIBUTE10 (PLBPPCS0TATTRIBUTE_IN[10], PLBPPCS0TATTRIBUTE[10]);
buf B_PLBPPCS0TATTRIBUTE11 (PLBPPCS0TATTRIBUTE_IN[11], PLBPPCS0TATTRIBUTE[11]);
buf B_PLBPPCS0TATTRIBUTE12 (PLBPPCS0TATTRIBUTE_IN[12], PLBPPCS0TATTRIBUTE[12]);
buf B_PLBPPCS0TATTRIBUTE13 (PLBPPCS0TATTRIBUTE_IN[13], PLBPPCS0TATTRIBUTE[13]);
buf B_PLBPPCS0TATTRIBUTE14 (PLBPPCS0TATTRIBUTE_IN[14], PLBPPCS0TATTRIBUTE[14]);
buf B_PLBPPCS0TATTRIBUTE15 (PLBPPCS0TATTRIBUTE_IN[15], PLBPPCS0TATTRIBUTE[15]);
buf B_PLBPPCS0TYPE0 (PLBPPCS0TYPE_IN[0], PLBPPCS0TYPE[0]);
buf B_PLBPPCS0TYPE1 (PLBPPCS0TYPE_IN[1], PLBPPCS0TYPE[1]);
buf B_PLBPPCS0TYPE2 (PLBPPCS0TYPE_IN[2], PLBPPCS0TYPE[2]);
buf B_PLBPPCS0UABUS28 (PLBPPCS0UABUS_IN[28], PLBPPCS0UABUS[28]);
buf B_PLBPPCS0UABUS29 (PLBPPCS0UABUS_IN[29], PLBPPCS0UABUS[29]);
buf B_PLBPPCS0UABUS30 (PLBPPCS0UABUS_IN[30], PLBPPCS0UABUS[30]);
buf B_PLBPPCS0UABUS31 (PLBPPCS0UABUS_IN[31], PLBPPCS0UABUS[31]);
buf B_PLBPPCS0WRBURST (PLBPPCS0WRBURST_IN, PLBPPCS0WRBURST);
buf B_PLBPPCS0WRDBUS0 (PLBPPCS0WRDBUS_IN[0], PLBPPCS0WRDBUS[0]);
buf B_PLBPPCS0WRDBUS1 (PLBPPCS0WRDBUS_IN[1], PLBPPCS0WRDBUS[1]);
buf B_PLBPPCS0WRDBUS2 (PLBPPCS0WRDBUS_IN[2], PLBPPCS0WRDBUS[2]);
buf B_PLBPPCS0WRDBUS3 (PLBPPCS0WRDBUS_IN[3], PLBPPCS0WRDBUS[3]);
buf B_PLBPPCS0WRDBUS4 (PLBPPCS0WRDBUS_IN[4], PLBPPCS0WRDBUS[4]);
buf B_PLBPPCS0WRDBUS5 (PLBPPCS0WRDBUS_IN[5], PLBPPCS0WRDBUS[5]);
buf B_PLBPPCS0WRDBUS6 (PLBPPCS0WRDBUS_IN[6], PLBPPCS0WRDBUS[6]);
buf B_PLBPPCS0WRDBUS7 (PLBPPCS0WRDBUS_IN[7], PLBPPCS0WRDBUS[7]);
buf B_PLBPPCS0WRDBUS8 (PLBPPCS0WRDBUS_IN[8], PLBPPCS0WRDBUS[8]);
buf B_PLBPPCS0WRDBUS9 (PLBPPCS0WRDBUS_IN[9], PLBPPCS0WRDBUS[9]);
buf B_PLBPPCS0WRDBUS10 (PLBPPCS0WRDBUS_IN[10], PLBPPCS0WRDBUS[10]);
buf B_PLBPPCS0WRDBUS11 (PLBPPCS0WRDBUS_IN[11], PLBPPCS0WRDBUS[11]);
buf B_PLBPPCS0WRDBUS12 (PLBPPCS0WRDBUS_IN[12], PLBPPCS0WRDBUS[12]);
buf B_PLBPPCS0WRDBUS13 (PLBPPCS0WRDBUS_IN[13], PLBPPCS0WRDBUS[13]);
buf B_PLBPPCS0WRDBUS14 (PLBPPCS0WRDBUS_IN[14], PLBPPCS0WRDBUS[14]);
buf B_PLBPPCS0WRDBUS15 (PLBPPCS0WRDBUS_IN[15], PLBPPCS0WRDBUS[15]);
buf B_PLBPPCS0WRDBUS16 (PLBPPCS0WRDBUS_IN[16], PLBPPCS0WRDBUS[16]);
buf B_PLBPPCS0WRDBUS17 (PLBPPCS0WRDBUS_IN[17], PLBPPCS0WRDBUS[17]);
buf B_PLBPPCS0WRDBUS18 (PLBPPCS0WRDBUS_IN[18], PLBPPCS0WRDBUS[18]);
buf B_PLBPPCS0WRDBUS19 (PLBPPCS0WRDBUS_IN[19], PLBPPCS0WRDBUS[19]);
buf B_PLBPPCS0WRDBUS20 (PLBPPCS0WRDBUS_IN[20], PLBPPCS0WRDBUS[20]);
buf B_PLBPPCS0WRDBUS21 (PLBPPCS0WRDBUS_IN[21], PLBPPCS0WRDBUS[21]);
buf B_PLBPPCS0WRDBUS22 (PLBPPCS0WRDBUS_IN[22], PLBPPCS0WRDBUS[22]);
buf B_PLBPPCS0WRDBUS23 (PLBPPCS0WRDBUS_IN[23], PLBPPCS0WRDBUS[23]);
buf B_PLBPPCS0WRDBUS24 (PLBPPCS0WRDBUS_IN[24], PLBPPCS0WRDBUS[24]);
buf B_PLBPPCS0WRDBUS25 (PLBPPCS0WRDBUS_IN[25], PLBPPCS0WRDBUS[25]);
buf B_PLBPPCS0WRDBUS26 (PLBPPCS0WRDBUS_IN[26], PLBPPCS0WRDBUS[26]);
buf B_PLBPPCS0WRDBUS27 (PLBPPCS0WRDBUS_IN[27], PLBPPCS0WRDBUS[27]);
buf B_PLBPPCS0WRDBUS28 (PLBPPCS0WRDBUS_IN[28], PLBPPCS0WRDBUS[28]);
buf B_PLBPPCS0WRDBUS29 (PLBPPCS0WRDBUS_IN[29], PLBPPCS0WRDBUS[29]);
buf B_PLBPPCS0WRDBUS30 (PLBPPCS0WRDBUS_IN[30], PLBPPCS0WRDBUS[30]);
buf B_PLBPPCS0WRDBUS31 (PLBPPCS0WRDBUS_IN[31], PLBPPCS0WRDBUS[31]);
buf B_PLBPPCS0WRDBUS32 (PLBPPCS0WRDBUS_IN[32], PLBPPCS0WRDBUS[32]);
buf B_PLBPPCS0WRDBUS33 (PLBPPCS0WRDBUS_IN[33], PLBPPCS0WRDBUS[33]);
buf B_PLBPPCS0WRDBUS34 (PLBPPCS0WRDBUS_IN[34], PLBPPCS0WRDBUS[34]);
buf B_PLBPPCS0WRDBUS35 (PLBPPCS0WRDBUS_IN[35], PLBPPCS0WRDBUS[35]);
buf B_PLBPPCS0WRDBUS36 (PLBPPCS0WRDBUS_IN[36], PLBPPCS0WRDBUS[36]);
buf B_PLBPPCS0WRDBUS37 (PLBPPCS0WRDBUS_IN[37], PLBPPCS0WRDBUS[37]);
buf B_PLBPPCS0WRDBUS38 (PLBPPCS0WRDBUS_IN[38], PLBPPCS0WRDBUS[38]);
buf B_PLBPPCS0WRDBUS39 (PLBPPCS0WRDBUS_IN[39], PLBPPCS0WRDBUS[39]);
buf B_PLBPPCS0WRDBUS40 (PLBPPCS0WRDBUS_IN[40], PLBPPCS0WRDBUS[40]);
buf B_PLBPPCS0WRDBUS41 (PLBPPCS0WRDBUS_IN[41], PLBPPCS0WRDBUS[41]);
buf B_PLBPPCS0WRDBUS42 (PLBPPCS0WRDBUS_IN[42], PLBPPCS0WRDBUS[42]);
buf B_PLBPPCS0WRDBUS43 (PLBPPCS0WRDBUS_IN[43], PLBPPCS0WRDBUS[43]);
buf B_PLBPPCS0WRDBUS44 (PLBPPCS0WRDBUS_IN[44], PLBPPCS0WRDBUS[44]);
buf B_PLBPPCS0WRDBUS45 (PLBPPCS0WRDBUS_IN[45], PLBPPCS0WRDBUS[45]);
buf B_PLBPPCS0WRDBUS46 (PLBPPCS0WRDBUS_IN[46], PLBPPCS0WRDBUS[46]);
buf B_PLBPPCS0WRDBUS47 (PLBPPCS0WRDBUS_IN[47], PLBPPCS0WRDBUS[47]);
buf B_PLBPPCS0WRDBUS48 (PLBPPCS0WRDBUS_IN[48], PLBPPCS0WRDBUS[48]);
buf B_PLBPPCS0WRDBUS49 (PLBPPCS0WRDBUS_IN[49], PLBPPCS0WRDBUS[49]);
buf B_PLBPPCS0WRDBUS50 (PLBPPCS0WRDBUS_IN[50], PLBPPCS0WRDBUS[50]);
buf B_PLBPPCS0WRDBUS51 (PLBPPCS0WRDBUS_IN[51], PLBPPCS0WRDBUS[51]);
buf B_PLBPPCS0WRDBUS52 (PLBPPCS0WRDBUS_IN[52], PLBPPCS0WRDBUS[52]);
buf B_PLBPPCS0WRDBUS53 (PLBPPCS0WRDBUS_IN[53], PLBPPCS0WRDBUS[53]);
buf B_PLBPPCS0WRDBUS54 (PLBPPCS0WRDBUS_IN[54], PLBPPCS0WRDBUS[54]);
buf B_PLBPPCS0WRDBUS55 (PLBPPCS0WRDBUS_IN[55], PLBPPCS0WRDBUS[55]);
buf B_PLBPPCS0WRDBUS56 (PLBPPCS0WRDBUS_IN[56], PLBPPCS0WRDBUS[56]);
buf B_PLBPPCS0WRDBUS57 (PLBPPCS0WRDBUS_IN[57], PLBPPCS0WRDBUS[57]);
buf B_PLBPPCS0WRDBUS58 (PLBPPCS0WRDBUS_IN[58], PLBPPCS0WRDBUS[58]);
buf B_PLBPPCS0WRDBUS59 (PLBPPCS0WRDBUS_IN[59], PLBPPCS0WRDBUS[59]);
buf B_PLBPPCS0WRDBUS60 (PLBPPCS0WRDBUS_IN[60], PLBPPCS0WRDBUS[60]);
buf B_PLBPPCS0WRDBUS61 (PLBPPCS0WRDBUS_IN[61], PLBPPCS0WRDBUS[61]);
buf B_PLBPPCS0WRDBUS62 (PLBPPCS0WRDBUS_IN[62], PLBPPCS0WRDBUS[62]);
buf B_PLBPPCS0WRDBUS63 (PLBPPCS0WRDBUS_IN[63], PLBPPCS0WRDBUS[63]);
buf B_PLBPPCS0WRDBUS64 (PLBPPCS0WRDBUS_IN[64], PLBPPCS0WRDBUS[64]);
buf B_PLBPPCS0WRDBUS65 (PLBPPCS0WRDBUS_IN[65], PLBPPCS0WRDBUS[65]);
buf B_PLBPPCS0WRDBUS66 (PLBPPCS0WRDBUS_IN[66], PLBPPCS0WRDBUS[66]);
buf B_PLBPPCS0WRDBUS67 (PLBPPCS0WRDBUS_IN[67], PLBPPCS0WRDBUS[67]);
buf B_PLBPPCS0WRDBUS68 (PLBPPCS0WRDBUS_IN[68], PLBPPCS0WRDBUS[68]);
buf B_PLBPPCS0WRDBUS69 (PLBPPCS0WRDBUS_IN[69], PLBPPCS0WRDBUS[69]);
buf B_PLBPPCS0WRDBUS70 (PLBPPCS0WRDBUS_IN[70], PLBPPCS0WRDBUS[70]);
buf B_PLBPPCS0WRDBUS71 (PLBPPCS0WRDBUS_IN[71], PLBPPCS0WRDBUS[71]);
buf B_PLBPPCS0WRDBUS72 (PLBPPCS0WRDBUS_IN[72], PLBPPCS0WRDBUS[72]);
buf B_PLBPPCS0WRDBUS73 (PLBPPCS0WRDBUS_IN[73], PLBPPCS0WRDBUS[73]);
buf B_PLBPPCS0WRDBUS74 (PLBPPCS0WRDBUS_IN[74], PLBPPCS0WRDBUS[74]);
buf B_PLBPPCS0WRDBUS75 (PLBPPCS0WRDBUS_IN[75], PLBPPCS0WRDBUS[75]);
buf B_PLBPPCS0WRDBUS76 (PLBPPCS0WRDBUS_IN[76], PLBPPCS0WRDBUS[76]);
buf B_PLBPPCS0WRDBUS77 (PLBPPCS0WRDBUS_IN[77], PLBPPCS0WRDBUS[77]);
buf B_PLBPPCS0WRDBUS78 (PLBPPCS0WRDBUS_IN[78], PLBPPCS0WRDBUS[78]);
buf B_PLBPPCS0WRDBUS79 (PLBPPCS0WRDBUS_IN[79], PLBPPCS0WRDBUS[79]);
buf B_PLBPPCS0WRDBUS80 (PLBPPCS0WRDBUS_IN[80], PLBPPCS0WRDBUS[80]);
buf B_PLBPPCS0WRDBUS81 (PLBPPCS0WRDBUS_IN[81], PLBPPCS0WRDBUS[81]);
buf B_PLBPPCS0WRDBUS82 (PLBPPCS0WRDBUS_IN[82], PLBPPCS0WRDBUS[82]);
buf B_PLBPPCS0WRDBUS83 (PLBPPCS0WRDBUS_IN[83], PLBPPCS0WRDBUS[83]);
buf B_PLBPPCS0WRDBUS84 (PLBPPCS0WRDBUS_IN[84], PLBPPCS0WRDBUS[84]);
buf B_PLBPPCS0WRDBUS85 (PLBPPCS0WRDBUS_IN[85], PLBPPCS0WRDBUS[85]);
buf B_PLBPPCS0WRDBUS86 (PLBPPCS0WRDBUS_IN[86], PLBPPCS0WRDBUS[86]);
buf B_PLBPPCS0WRDBUS87 (PLBPPCS0WRDBUS_IN[87], PLBPPCS0WRDBUS[87]);
buf B_PLBPPCS0WRDBUS88 (PLBPPCS0WRDBUS_IN[88], PLBPPCS0WRDBUS[88]);
buf B_PLBPPCS0WRDBUS89 (PLBPPCS0WRDBUS_IN[89], PLBPPCS0WRDBUS[89]);
buf B_PLBPPCS0WRDBUS90 (PLBPPCS0WRDBUS_IN[90], PLBPPCS0WRDBUS[90]);
buf B_PLBPPCS0WRDBUS91 (PLBPPCS0WRDBUS_IN[91], PLBPPCS0WRDBUS[91]);
buf B_PLBPPCS0WRDBUS92 (PLBPPCS0WRDBUS_IN[92], PLBPPCS0WRDBUS[92]);
buf B_PLBPPCS0WRDBUS93 (PLBPPCS0WRDBUS_IN[93], PLBPPCS0WRDBUS[93]);
buf B_PLBPPCS0WRDBUS94 (PLBPPCS0WRDBUS_IN[94], PLBPPCS0WRDBUS[94]);
buf B_PLBPPCS0WRDBUS95 (PLBPPCS0WRDBUS_IN[95], PLBPPCS0WRDBUS[95]);
buf B_PLBPPCS0WRDBUS96 (PLBPPCS0WRDBUS_IN[96], PLBPPCS0WRDBUS[96]);
buf B_PLBPPCS0WRDBUS97 (PLBPPCS0WRDBUS_IN[97], PLBPPCS0WRDBUS[97]);
buf B_PLBPPCS0WRDBUS98 (PLBPPCS0WRDBUS_IN[98], PLBPPCS0WRDBUS[98]);
buf B_PLBPPCS0WRDBUS99 (PLBPPCS0WRDBUS_IN[99], PLBPPCS0WRDBUS[99]);
buf B_PLBPPCS0WRDBUS100 (PLBPPCS0WRDBUS_IN[100], PLBPPCS0WRDBUS[100]);
buf B_PLBPPCS0WRDBUS101 (PLBPPCS0WRDBUS_IN[101], PLBPPCS0WRDBUS[101]);
buf B_PLBPPCS0WRDBUS102 (PLBPPCS0WRDBUS_IN[102], PLBPPCS0WRDBUS[102]);
buf B_PLBPPCS0WRDBUS103 (PLBPPCS0WRDBUS_IN[103], PLBPPCS0WRDBUS[103]);
buf B_PLBPPCS0WRDBUS104 (PLBPPCS0WRDBUS_IN[104], PLBPPCS0WRDBUS[104]);
buf B_PLBPPCS0WRDBUS105 (PLBPPCS0WRDBUS_IN[105], PLBPPCS0WRDBUS[105]);
buf B_PLBPPCS0WRDBUS106 (PLBPPCS0WRDBUS_IN[106], PLBPPCS0WRDBUS[106]);
buf B_PLBPPCS0WRDBUS107 (PLBPPCS0WRDBUS_IN[107], PLBPPCS0WRDBUS[107]);
buf B_PLBPPCS0WRDBUS108 (PLBPPCS0WRDBUS_IN[108], PLBPPCS0WRDBUS[108]);
buf B_PLBPPCS0WRDBUS109 (PLBPPCS0WRDBUS_IN[109], PLBPPCS0WRDBUS[109]);
buf B_PLBPPCS0WRDBUS110 (PLBPPCS0WRDBUS_IN[110], PLBPPCS0WRDBUS[110]);
buf B_PLBPPCS0WRDBUS111 (PLBPPCS0WRDBUS_IN[111], PLBPPCS0WRDBUS[111]);
buf B_PLBPPCS0WRDBUS112 (PLBPPCS0WRDBUS_IN[112], PLBPPCS0WRDBUS[112]);
buf B_PLBPPCS0WRDBUS113 (PLBPPCS0WRDBUS_IN[113], PLBPPCS0WRDBUS[113]);
buf B_PLBPPCS0WRDBUS114 (PLBPPCS0WRDBUS_IN[114], PLBPPCS0WRDBUS[114]);
buf B_PLBPPCS0WRDBUS115 (PLBPPCS0WRDBUS_IN[115], PLBPPCS0WRDBUS[115]);
buf B_PLBPPCS0WRDBUS116 (PLBPPCS0WRDBUS_IN[116], PLBPPCS0WRDBUS[116]);
buf B_PLBPPCS0WRDBUS117 (PLBPPCS0WRDBUS_IN[117], PLBPPCS0WRDBUS[117]);
buf B_PLBPPCS0WRDBUS118 (PLBPPCS0WRDBUS_IN[118], PLBPPCS0WRDBUS[118]);
buf B_PLBPPCS0WRDBUS119 (PLBPPCS0WRDBUS_IN[119], PLBPPCS0WRDBUS[119]);
buf B_PLBPPCS0WRDBUS120 (PLBPPCS0WRDBUS_IN[120], PLBPPCS0WRDBUS[120]);
buf B_PLBPPCS0WRDBUS121 (PLBPPCS0WRDBUS_IN[121], PLBPPCS0WRDBUS[121]);
buf B_PLBPPCS0WRDBUS122 (PLBPPCS0WRDBUS_IN[122], PLBPPCS0WRDBUS[122]);
buf B_PLBPPCS0WRDBUS123 (PLBPPCS0WRDBUS_IN[123], PLBPPCS0WRDBUS[123]);
buf B_PLBPPCS0WRDBUS124 (PLBPPCS0WRDBUS_IN[124], PLBPPCS0WRDBUS[124]);
buf B_PLBPPCS0WRDBUS125 (PLBPPCS0WRDBUS_IN[125], PLBPPCS0WRDBUS[125]);
buf B_PLBPPCS0WRDBUS126 (PLBPPCS0WRDBUS_IN[126], PLBPPCS0WRDBUS[126]);
buf B_PLBPPCS0WRDBUS127 (PLBPPCS0WRDBUS_IN[127], PLBPPCS0WRDBUS[127]);
buf B_PLBPPCS0WRPENDPRI0 (PLBPPCS0WRPENDPRI_IN[0], PLBPPCS0WRPENDPRI[0]);
buf B_PLBPPCS0WRPENDPRI1 (PLBPPCS0WRPENDPRI_IN[1], PLBPPCS0WRPENDPRI[1]);
buf B_PLBPPCS0WRPENDREQ (PLBPPCS0WRPENDREQ_IN, PLBPPCS0WRPENDREQ);
buf B_PLBPPCS0WRPRIM (PLBPPCS0WRPRIM_IN, PLBPPCS0WRPRIM);
buf B_PLBPPCS1ABORT (PLBPPCS1ABORT_IN, PLBPPCS1ABORT);
buf B_PLBPPCS1ABUS0 (PLBPPCS1ABUS_IN[0], PLBPPCS1ABUS[0]);
buf B_PLBPPCS1ABUS1 (PLBPPCS1ABUS_IN[1], PLBPPCS1ABUS[1]);
buf B_PLBPPCS1ABUS2 (PLBPPCS1ABUS_IN[2], PLBPPCS1ABUS[2]);
buf B_PLBPPCS1ABUS3 (PLBPPCS1ABUS_IN[3], PLBPPCS1ABUS[3]);
buf B_PLBPPCS1ABUS4 (PLBPPCS1ABUS_IN[4], PLBPPCS1ABUS[4]);
buf B_PLBPPCS1ABUS5 (PLBPPCS1ABUS_IN[5], PLBPPCS1ABUS[5]);
buf B_PLBPPCS1ABUS6 (PLBPPCS1ABUS_IN[6], PLBPPCS1ABUS[6]);
buf B_PLBPPCS1ABUS7 (PLBPPCS1ABUS_IN[7], PLBPPCS1ABUS[7]);
buf B_PLBPPCS1ABUS8 (PLBPPCS1ABUS_IN[8], PLBPPCS1ABUS[8]);
buf B_PLBPPCS1ABUS9 (PLBPPCS1ABUS_IN[9], PLBPPCS1ABUS[9]);
buf B_PLBPPCS1ABUS10 (PLBPPCS1ABUS_IN[10], PLBPPCS1ABUS[10]);
buf B_PLBPPCS1ABUS11 (PLBPPCS1ABUS_IN[11], PLBPPCS1ABUS[11]);
buf B_PLBPPCS1ABUS12 (PLBPPCS1ABUS_IN[12], PLBPPCS1ABUS[12]);
buf B_PLBPPCS1ABUS13 (PLBPPCS1ABUS_IN[13], PLBPPCS1ABUS[13]);
buf B_PLBPPCS1ABUS14 (PLBPPCS1ABUS_IN[14], PLBPPCS1ABUS[14]);
buf B_PLBPPCS1ABUS15 (PLBPPCS1ABUS_IN[15], PLBPPCS1ABUS[15]);
buf B_PLBPPCS1ABUS16 (PLBPPCS1ABUS_IN[16], PLBPPCS1ABUS[16]);
buf B_PLBPPCS1ABUS17 (PLBPPCS1ABUS_IN[17], PLBPPCS1ABUS[17]);
buf B_PLBPPCS1ABUS18 (PLBPPCS1ABUS_IN[18], PLBPPCS1ABUS[18]);
buf B_PLBPPCS1ABUS19 (PLBPPCS1ABUS_IN[19], PLBPPCS1ABUS[19]);
buf B_PLBPPCS1ABUS20 (PLBPPCS1ABUS_IN[20], PLBPPCS1ABUS[20]);
buf B_PLBPPCS1ABUS21 (PLBPPCS1ABUS_IN[21], PLBPPCS1ABUS[21]);
buf B_PLBPPCS1ABUS22 (PLBPPCS1ABUS_IN[22], PLBPPCS1ABUS[22]);
buf B_PLBPPCS1ABUS23 (PLBPPCS1ABUS_IN[23], PLBPPCS1ABUS[23]);
buf B_PLBPPCS1ABUS24 (PLBPPCS1ABUS_IN[24], PLBPPCS1ABUS[24]);
buf B_PLBPPCS1ABUS25 (PLBPPCS1ABUS_IN[25], PLBPPCS1ABUS[25]);
buf B_PLBPPCS1ABUS26 (PLBPPCS1ABUS_IN[26], PLBPPCS1ABUS[26]);
buf B_PLBPPCS1ABUS27 (PLBPPCS1ABUS_IN[27], PLBPPCS1ABUS[27]);
buf B_PLBPPCS1ABUS28 (PLBPPCS1ABUS_IN[28], PLBPPCS1ABUS[28]);
buf B_PLBPPCS1ABUS29 (PLBPPCS1ABUS_IN[29], PLBPPCS1ABUS[29]);
buf B_PLBPPCS1ABUS30 (PLBPPCS1ABUS_IN[30], PLBPPCS1ABUS[30]);
buf B_PLBPPCS1ABUS31 (PLBPPCS1ABUS_IN[31], PLBPPCS1ABUS[31]);
buf B_PLBPPCS1BE0 (PLBPPCS1BE_IN[0], PLBPPCS1BE[0]);
buf B_PLBPPCS1BE1 (PLBPPCS1BE_IN[1], PLBPPCS1BE[1]);
buf B_PLBPPCS1BE2 (PLBPPCS1BE_IN[2], PLBPPCS1BE[2]);
buf B_PLBPPCS1BE3 (PLBPPCS1BE_IN[3], PLBPPCS1BE[3]);
buf B_PLBPPCS1BE4 (PLBPPCS1BE_IN[4], PLBPPCS1BE[4]);
buf B_PLBPPCS1BE5 (PLBPPCS1BE_IN[5], PLBPPCS1BE[5]);
buf B_PLBPPCS1BE6 (PLBPPCS1BE_IN[6], PLBPPCS1BE[6]);
buf B_PLBPPCS1BE7 (PLBPPCS1BE_IN[7], PLBPPCS1BE[7]);
buf B_PLBPPCS1BE8 (PLBPPCS1BE_IN[8], PLBPPCS1BE[8]);
buf B_PLBPPCS1BE9 (PLBPPCS1BE_IN[9], PLBPPCS1BE[9]);
buf B_PLBPPCS1BE10 (PLBPPCS1BE_IN[10], PLBPPCS1BE[10]);
buf B_PLBPPCS1BE11 (PLBPPCS1BE_IN[11], PLBPPCS1BE[11]);
buf B_PLBPPCS1BE12 (PLBPPCS1BE_IN[12], PLBPPCS1BE[12]);
buf B_PLBPPCS1BE13 (PLBPPCS1BE_IN[13], PLBPPCS1BE[13]);
buf B_PLBPPCS1BE14 (PLBPPCS1BE_IN[14], PLBPPCS1BE[14]);
buf B_PLBPPCS1BE15 (PLBPPCS1BE_IN[15], PLBPPCS1BE[15]);
buf B_PLBPPCS1BUSLOCK (PLBPPCS1BUSLOCK_IN, PLBPPCS1BUSLOCK);
buf B_PLBPPCS1LOCKERR (PLBPPCS1LOCKERR_IN, PLBPPCS1LOCKERR);
buf B_PLBPPCS1MASTERID0 (PLBPPCS1MASTERID_IN[0], PLBPPCS1MASTERID[0]);
buf B_PLBPPCS1MASTERID1 (PLBPPCS1MASTERID_IN[1], PLBPPCS1MASTERID[1]);
buf B_PLBPPCS1MSIZE0 (PLBPPCS1MSIZE_IN[0], PLBPPCS1MSIZE[0]);
buf B_PLBPPCS1MSIZE1 (PLBPPCS1MSIZE_IN[1], PLBPPCS1MSIZE[1]);
buf B_PLBPPCS1PAVALID (PLBPPCS1PAVALID_IN, PLBPPCS1PAVALID);
buf B_PLBPPCS1RDBURST (PLBPPCS1RDBURST_IN, PLBPPCS1RDBURST);
buf B_PLBPPCS1RDPENDPRI0 (PLBPPCS1RDPENDPRI_IN[0], PLBPPCS1RDPENDPRI[0]);
buf B_PLBPPCS1RDPENDPRI1 (PLBPPCS1RDPENDPRI_IN[1], PLBPPCS1RDPENDPRI[1]);
buf B_PLBPPCS1RDPENDREQ (PLBPPCS1RDPENDREQ_IN, PLBPPCS1RDPENDREQ);
buf B_PLBPPCS1RDPRIM (PLBPPCS1RDPRIM_IN, PLBPPCS1RDPRIM);
buf B_PLBPPCS1REQPRI0 (PLBPPCS1REQPRI_IN[0], PLBPPCS1REQPRI[0]);
buf B_PLBPPCS1REQPRI1 (PLBPPCS1REQPRI_IN[1], PLBPPCS1REQPRI[1]);
buf B_PLBPPCS1SAVALID (PLBPPCS1SAVALID_IN, PLBPPCS1SAVALID);
buf B_PLBPPCS1SIZE0 (PLBPPCS1SIZE_IN[0], PLBPPCS1SIZE[0]);
buf B_PLBPPCS1SIZE1 (PLBPPCS1SIZE_IN[1], PLBPPCS1SIZE[1]);
buf B_PLBPPCS1SIZE2 (PLBPPCS1SIZE_IN[2], PLBPPCS1SIZE[2]);
buf B_PLBPPCS1SIZE3 (PLBPPCS1SIZE_IN[3], PLBPPCS1SIZE[3]);
buf B_PLBPPCS1TATTRIBUTE0 (PLBPPCS1TATTRIBUTE_IN[0], PLBPPCS1TATTRIBUTE[0]);
buf B_PLBPPCS1TATTRIBUTE1 (PLBPPCS1TATTRIBUTE_IN[1], PLBPPCS1TATTRIBUTE[1]);
buf B_PLBPPCS1TATTRIBUTE2 (PLBPPCS1TATTRIBUTE_IN[2], PLBPPCS1TATTRIBUTE[2]);
buf B_PLBPPCS1TATTRIBUTE3 (PLBPPCS1TATTRIBUTE_IN[3], PLBPPCS1TATTRIBUTE[3]);
buf B_PLBPPCS1TATTRIBUTE4 (PLBPPCS1TATTRIBUTE_IN[4], PLBPPCS1TATTRIBUTE[4]);
buf B_PLBPPCS1TATTRIBUTE5 (PLBPPCS1TATTRIBUTE_IN[5], PLBPPCS1TATTRIBUTE[5]);
buf B_PLBPPCS1TATTRIBUTE6 (PLBPPCS1TATTRIBUTE_IN[6], PLBPPCS1TATTRIBUTE[6]);
buf B_PLBPPCS1TATTRIBUTE7 (PLBPPCS1TATTRIBUTE_IN[7], PLBPPCS1TATTRIBUTE[7]);
buf B_PLBPPCS1TATTRIBUTE8 (PLBPPCS1TATTRIBUTE_IN[8], PLBPPCS1TATTRIBUTE[8]);
buf B_PLBPPCS1TATTRIBUTE9 (PLBPPCS1TATTRIBUTE_IN[9], PLBPPCS1TATTRIBUTE[9]);
buf B_PLBPPCS1TATTRIBUTE10 (PLBPPCS1TATTRIBUTE_IN[10], PLBPPCS1TATTRIBUTE[10]);
buf B_PLBPPCS1TATTRIBUTE11 (PLBPPCS1TATTRIBUTE_IN[11], PLBPPCS1TATTRIBUTE[11]);
buf B_PLBPPCS1TATTRIBUTE12 (PLBPPCS1TATTRIBUTE_IN[12], PLBPPCS1TATTRIBUTE[12]);
buf B_PLBPPCS1TATTRIBUTE13 (PLBPPCS1TATTRIBUTE_IN[13], PLBPPCS1TATTRIBUTE[13]);
buf B_PLBPPCS1TATTRIBUTE14 (PLBPPCS1TATTRIBUTE_IN[14], PLBPPCS1TATTRIBUTE[14]);
buf B_PLBPPCS1TATTRIBUTE15 (PLBPPCS1TATTRIBUTE_IN[15], PLBPPCS1TATTRIBUTE[15]);
buf B_PLBPPCS1TYPE0 (PLBPPCS1TYPE_IN[0], PLBPPCS1TYPE[0]);
buf B_PLBPPCS1TYPE1 (PLBPPCS1TYPE_IN[1], PLBPPCS1TYPE[1]);
buf B_PLBPPCS1TYPE2 (PLBPPCS1TYPE_IN[2], PLBPPCS1TYPE[2]);
buf B_PLBPPCS1UABUS28 (PLBPPCS1UABUS_IN[28], PLBPPCS1UABUS[28]);
buf B_PLBPPCS1UABUS29 (PLBPPCS1UABUS_IN[29], PLBPPCS1UABUS[29]);
buf B_PLBPPCS1UABUS30 (PLBPPCS1UABUS_IN[30], PLBPPCS1UABUS[30]);
buf B_PLBPPCS1UABUS31 (PLBPPCS1UABUS_IN[31], PLBPPCS1UABUS[31]);
buf B_PLBPPCS1WRBURST (PLBPPCS1WRBURST_IN, PLBPPCS1WRBURST);
buf B_PLBPPCS1WRDBUS0 (PLBPPCS1WRDBUS_IN[0], PLBPPCS1WRDBUS[0]);
buf B_PLBPPCS1WRDBUS1 (PLBPPCS1WRDBUS_IN[1], PLBPPCS1WRDBUS[1]);
buf B_PLBPPCS1WRDBUS2 (PLBPPCS1WRDBUS_IN[2], PLBPPCS1WRDBUS[2]);
buf B_PLBPPCS1WRDBUS3 (PLBPPCS1WRDBUS_IN[3], PLBPPCS1WRDBUS[3]);
buf B_PLBPPCS1WRDBUS4 (PLBPPCS1WRDBUS_IN[4], PLBPPCS1WRDBUS[4]);
buf B_PLBPPCS1WRDBUS5 (PLBPPCS1WRDBUS_IN[5], PLBPPCS1WRDBUS[5]);
buf B_PLBPPCS1WRDBUS6 (PLBPPCS1WRDBUS_IN[6], PLBPPCS1WRDBUS[6]);
buf B_PLBPPCS1WRDBUS7 (PLBPPCS1WRDBUS_IN[7], PLBPPCS1WRDBUS[7]);
buf B_PLBPPCS1WRDBUS8 (PLBPPCS1WRDBUS_IN[8], PLBPPCS1WRDBUS[8]);
buf B_PLBPPCS1WRDBUS9 (PLBPPCS1WRDBUS_IN[9], PLBPPCS1WRDBUS[9]);
buf B_PLBPPCS1WRDBUS10 (PLBPPCS1WRDBUS_IN[10], PLBPPCS1WRDBUS[10]);
buf B_PLBPPCS1WRDBUS11 (PLBPPCS1WRDBUS_IN[11], PLBPPCS1WRDBUS[11]);
buf B_PLBPPCS1WRDBUS12 (PLBPPCS1WRDBUS_IN[12], PLBPPCS1WRDBUS[12]);
buf B_PLBPPCS1WRDBUS13 (PLBPPCS1WRDBUS_IN[13], PLBPPCS1WRDBUS[13]);
buf B_PLBPPCS1WRDBUS14 (PLBPPCS1WRDBUS_IN[14], PLBPPCS1WRDBUS[14]);
buf B_PLBPPCS1WRDBUS15 (PLBPPCS1WRDBUS_IN[15], PLBPPCS1WRDBUS[15]);
buf B_PLBPPCS1WRDBUS16 (PLBPPCS1WRDBUS_IN[16], PLBPPCS1WRDBUS[16]);
buf B_PLBPPCS1WRDBUS17 (PLBPPCS1WRDBUS_IN[17], PLBPPCS1WRDBUS[17]);
buf B_PLBPPCS1WRDBUS18 (PLBPPCS1WRDBUS_IN[18], PLBPPCS1WRDBUS[18]);
buf B_PLBPPCS1WRDBUS19 (PLBPPCS1WRDBUS_IN[19], PLBPPCS1WRDBUS[19]);
buf B_PLBPPCS1WRDBUS20 (PLBPPCS1WRDBUS_IN[20], PLBPPCS1WRDBUS[20]);
buf B_PLBPPCS1WRDBUS21 (PLBPPCS1WRDBUS_IN[21], PLBPPCS1WRDBUS[21]);
buf B_PLBPPCS1WRDBUS22 (PLBPPCS1WRDBUS_IN[22], PLBPPCS1WRDBUS[22]);
buf B_PLBPPCS1WRDBUS23 (PLBPPCS1WRDBUS_IN[23], PLBPPCS1WRDBUS[23]);
buf B_PLBPPCS1WRDBUS24 (PLBPPCS1WRDBUS_IN[24], PLBPPCS1WRDBUS[24]);
buf B_PLBPPCS1WRDBUS25 (PLBPPCS1WRDBUS_IN[25], PLBPPCS1WRDBUS[25]);
buf B_PLBPPCS1WRDBUS26 (PLBPPCS1WRDBUS_IN[26], PLBPPCS1WRDBUS[26]);
buf B_PLBPPCS1WRDBUS27 (PLBPPCS1WRDBUS_IN[27], PLBPPCS1WRDBUS[27]);
buf B_PLBPPCS1WRDBUS28 (PLBPPCS1WRDBUS_IN[28], PLBPPCS1WRDBUS[28]);
buf B_PLBPPCS1WRDBUS29 (PLBPPCS1WRDBUS_IN[29], PLBPPCS1WRDBUS[29]);
buf B_PLBPPCS1WRDBUS30 (PLBPPCS1WRDBUS_IN[30], PLBPPCS1WRDBUS[30]);
buf B_PLBPPCS1WRDBUS31 (PLBPPCS1WRDBUS_IN[31], PLBPPCS1WRDBUS[31]);
buf B_PLBPPCS1WRDBUS32 (PLBPPCS1WRDBUS_IN[32], PLBPPCS1WRDBUS[32]);
buf B_PLBPPCS1WRDBUS33 (PLBPPCS1WRDBUS_IN[33], PLBPPCS1WRDBUS[33]);
buf B_PLBPPCS1WRDBUS34 (PLBPPCS1WRDBUS_IN[34], PLBPPCS1WRDBUS[34]);
buf B_PLBPPCS1WRDBUS35 (PLBPPCS1WRDBUS_IN[35], PLBPPCS1WRDBUS[35]);
buf B_PLBPPCS1WRDBUS36 (PLBPPCS1WRDBUS_IN[36], PLBPPCS1WRDBUS[36]);
buf B_PLBPPCS1WRDBUS37 (PLBPPCS1WRDBUS_IN[37], PLBPPCS1WRDBUS[37]);
buf B_PLBPPCS1WRDBUS38 (PLBPPCS1WRDBUS_IN[38], PLBPPCS1WRDBUS[38]);
buf B_PLBPPCS1WRDBUS39 (PLBPPCS1WRDBUS_IN[39], PLBPPCS1WRDBUS[39]);
buf B_PLBPPCS1WRDBUS40 (PLBPPCS1WRDBUS_IN[40], PLBPPCS1WRDBUS[40]);
buf B_PLBPPCS1WRDBUS41 (PLBPPCS1WRDBUS_IN[41], PLBPPCS1WRDBUS[41]);
buf B_PLBPPCS1WRDBUS42 (PLBPPCS1WRDBUS_IN[42], PLBPPCS1WRDBUS[42]);
buf B_PLBPPCS1WRDBUS43 (PLBPPCS1WRDBUS_IN[43], PLBPPCS1WRDBUS[43]);
buf B_PLBPPCS1WRDBUS44 (PLBPPCS1WRDBUS_IN[44], PLBPPCS1WRDBUS[44]);
buf B_PLBPPCS1WRDBUS45 (PLBPPCS1WRDBUS_IN[45], PLBPPCS1WRDBUS[45]);
buf B_PLBPPCS1WRDBUS46 (PLBPPCS1WRDBUS_IN[46], PLBPPCS1WRDBUS[46]);
buf B_PLBPPCS1WRDBUS47 (PLBPPCS1WRDBUS_IN[47], PLBPPCS1WRDBUS[47]);
buf B_PLBPPCS1WRDBUS48 (PLBPPCS1WRDBUS_IN[48], PLBPPCS1WRDBUS[48]);
buf B_PLBPPCS1WRDBUS49 (PLBPPCS1WRDBUS_IN[49], PLBPPCS1WRDBUS[49]);
buf B_PLBPPCS1WRDBUS50 (PLBPPCS1WRDBUS_IN[50], PLBPPCS1WRDBUS[50]);
buf B_PLBPPCS1WRDBUS51 (PLBPPCS1WRDBUS_IN[51], PLBPPCS1WRDBUS[51]);
buf B_PLBPPCS1WRDBUS52 (PLBPPCS1WRDBUS_IN[52], PLBPPCS1WRDBUS[52]);
buf B_PLBPPCS1WRDBUS53 (PLBPPCS1WRDBUS_IN[53], PLBPPCS1WRDBUS[53]);
buf B_PLBPPCS1WRDBUS54 (PLBPPCS1WRDBUS_IN[54], PLBPPCS1WRDBUS[54]);
buf B_PLBPPCS1WRDBUS55 (PLBPPCS1WRDBUS_IN[55], PLBPPCS1WRDBUS[55]);
buf B_PLBPPCS1WRDBUS56 (PLBPPCS1WRDBUS_IN[56], PLBPPCS1WRDBUS[56]);
buf B_PLBPPCS1WRDBUS57 (PLBPPCS1WRDBUS_IN[57], PLBPPCS1WRDBUS[57]);
buf B_PLBPPCS1WRDBUS58 (PLBPPCS1WRDBUS_IN[58], PLBPPCS1WRDBUS[58]);
buf B_PLBPPCS1WRDBUS59 (PLBPPCS1WRDBUS_IN[59], PLBPPCS1WRDBUS[59]);
buf B_PLBPPCS1WRDBUS60 (PLBPPCS1WRDBUS_IN[60], PLBPPCS1WRDBUS[60]);
buf B_PLBPPCS1WRDBUS61 (PLBPPCS1WRDBUS_IN[61], PLBPPCS1WRDBUS[61]);
buf B_PLBPPCS1WRDBUS62 (PLBPPCS1WRDBUS_IN[62], PLBPPCS1WRDBUS[62]);
buf B_PLBPPCS1WRDBUS63 (PLBPPCS1WRDBUS_IN[63], PLBPPCS1WRDBUS[63]);
buf B_PLBPPCS1WRDBUS64 (PLBPPCS1WRDBUS_IN[64], PLBPPCS1WRDBUS[64]);
buf B_PLBPPCS1WRDBUS65 (PLBPPCS1WRDBUS_IN[65], PLBPPCS1WRDBUS[65]);
buf B_PLBPPCS1WRDBUS66 (PLBPPCS1WRDBUS_IN[66], PLBPPCS1WRDBUS[66]);
buf B_PLBPPCS1WRDBUS67 (PLBPPCS1WRDBUS_IN[67], PLBPPCS1WRDBUS[67]);
buf B_PLBPPCS1WRDBUS68 (PLBPPCS1WRDBUS_IN[68], PLBPPCS1WRDBUS[68]);
buf B_PLBPPCS1WRDBUS69 (PLBPPCS1WRDBUS_IN[69], PLBPPCS1WRDBUS[69]);
buf B_PLBPPCS1WRDBUS70 (PLBPPCS1WRDBUS_IN[70], PLBPPCS1WRDBUS[70]);
buf B_PLBPPCS1WRDBUS71 (PLBPPCS1WRDBUS_IN[71], PLBPPCS1WRDBUS[71]);
buf B_PLBPPCS1WRDBUS72 (PLBPPCS1WRDBUS_IN[72], PLBPPCS1WRDBUS[72]);
buf B_PLBPPCS1WRDBUS73 (PLBPPCS1WRDBUS_IN[73], PLBPPCS1WRDBUS[73]);
buf B_PLBPPCS1WRDBUS74 (PLBPPCS1WRDBUS_IN[74], PLBPPCS1WRDBUS[74]);
buf B_PLBPPCS1WRDBUS75 (PLBPPCS1WRDBUS_IN[75], PLBPPCS1WRDBUS[75]);
buf B_PLBPPCS1WRDBUS76 (PLBPPCS1WRDBUS_IN[76], PLBPPCS1WRDBUS[76]);
buf B_PLBPPCS1WRDBUS77 (PLBPPCS1WRDBUS_IN[77], PLBPPCS1WRDBUS[77]);
buf B_PLBPPCS1WRDBUS78 (PLBPPCS1WRDBUS_IN[78], PLBPPCS1WRDBUS[78]);
buf B_PLBPPCS1WRDBUS79 (PLBPPCS1WRDBUS_IN[79], PLBPPCS1WRDBUS[79]);
buf B_PLBPPCS1WRDBUS80 (PLBPPCS1WRDBUS_IN[80], PLBPPCS1WRDBUS[80]);
buf B_PLBPPCS1WRDBUS81 (PLBPPCS1WRDBUS_IN[81], PLBPPCS1WRDBUS[81]);
buf B_PLBPPCS1WRDBUS82 (PLBPPCS1WRDBUS_IN[82], PLBPPCS1WRDBUS[82]);
buf B_PLBPPCS1WRDBUS83 (PLBPPCS1WRDBUS_IN[83], PLBPPCS1WRDBUS[83]);
buf B_PLBPPCS1WRDBUS84 (PLBPPCS1WRDBUS_IN[84], PLBPPCS1WRDBUS[84]);
buf B_PLBPPCS1WRDBUS85 (PLBPPCS1WRDBUS_IN[85], PLBPPCS1WRDBUS[85]);
buf B_PLBPPCS1WRDBUS86 (PLBPPCS1WRDBUS_IN[86], PLBPPCS1WRDBUS[86]);
buf B_PLBPPCS1WRDBUS87 (PLBPPCS1WRDBUS_IN[87], PLBPPCS1WRDBUS[87]);
buf B_PLBPPCS1WRDBUS88 (PLBPPCS1WRDBUS_IN[88], PLBPPCS1WRDBUS[88]);
buf B_PLBPPCS1WRDBUS89 (PLBPPCS1WRDBUS_IN[89], PLBPPCS1WRDBUS[89]);
buf B_PLBPPCS1WRDBUS90 (PLBPPCS1WRDBUS_IN[90], PLBPPCS1WRDBUS[90]);
buf B_PLBPPCS1WRDBUS91 (PLBPPCS1WRDBUS_IN[91], PLBPPCS1WRDBUS[91]);
buf B_PLBPPCS1WRDBUS92 (PLBPPCS1WRDBUS_IN[92], PLBPPCS1WRDBUS[92]);
buf B_PLBPPCS1WRDBUS93 (PLBPPCS1WRDBUS_IN[93], PLBPPCS1WRDBUS[93]);
buf B_PLBPPCS1WRDBUS94 (PLBPPCS1WRDBUS_IN[94], PLBPPCS1WRDBUS[94]);
buf B_PLBPPCS1WRDBUS95 (PLBPPCS1WRDBUS_IN[95], PLBPPCS1WRDBUS[95]);
buf B_PLBPPCS1WRDBUS96 (PLBPPCS1WRDBUS_IN[96], PLBPPCS1WRDBUS[96]);
buf B_PLBPPCS1WRDBUS97 (PLBPPCS1WRDBUS_IN[97], PLBPPCS1WRDBUS[97]);
buf B_PLBPPCS1WRDBUS98 (PLBPPCS1WRDBUS_IN[98], PLBPPCS1WRDBUS[98]);
buf B_PLBPPCS1WRDBUS99 (PLBPPCS1WRDBUS_IN[99], PLBPPCS1WRDBUS[99]);
buf B_PLBPPCS1WRDBUS100 (PLBPPCS1WRDBUS_IN[100], PLBPPCS1WRDBUS[100]);
buf B_PLBPPCS1WRDBUS101 (PLBPPCS1WRDBUS_IN[101], PLBPPCS1WRDBUS[101]);
buf B_PLBPPCS1WRDBUS102 (PLBPPCS1WRDBUS_IN[102], PLBPPCS1WRDBUS[102]);
buf B_PLBPPCS1WRDBUS103 (PLBPPCS1WRDBUS_IN[103], PLBPPCS1WRDBUS[103]);
buf B_PLBPPCS1WRDBUS104 (PLBPPCS1WRDBUS_IN[104], PLBPPCS1WRDBUS[104]);
buf B_PLBPPCS1WRDBUS105 (PLBPPCS1WRDBUS_IN[105], PLBPPCS1WRDBUS[105]);
buf B_PLBPPCS1WRDBUS106 (PLBPPCS1WRDBUS_IN[106], PLBPPCS1WRDBUS[106]);
buf B_PLBPPCS1WRDBUS107 (PLBPPCS1WRDBUS_IN[107], PLBPPCS1WRDBUS[107]);
buf B_PLBPPCS1WRDBUS108 (PLBPPCS1WRDBUS_IN[108], PLBPPCS1WRDBUS[108]);
buf B_PLBPPCS1WRDBUS109 (PLBPPCS1WRDBUS_IN[109], PLBPPCS1WRDBUS[109]);
buf B_PLBPPCS1WRDBUS110 (PLBPPCS1WRDBUS_IN[110], PLBPPCS1WRDBUS[110]);
buf B_PLBPPCS1WRDBUS111 (PLBPPCS1WRDBUS_IN[111], PLBPPCS1WRDBUS[111]);
buf B_PLBPPCS1WRDBUS112 (PLBPPCS1WRDBUS_IN[112], PLBPPCS1WRDBUS[112]);
buf B_PLBPPCS1WRDBUS113 (PLBPPCS1WRDBUS_IN[113], PLBPPCS1WRDBUS[113]);
buf B_PLBPPCS1WRDBUS114 (PLBPPCS1WRDBUS_IN[114], PLBPPCS1WRDBUS[114]);
buf B_PLBPPCS1WRDBUS115 (PLBPPCS1WRDBUS_IN[115], PLBPPCS1WRDBUS[115]);
buf B_PLBPPCS1WRDBUS116 (PLBPPCS1WRDBUS_IN[116], PLBPPCS1WRDBUS[116]);
buf B_PLBPPCS1WRDBUS117 (PLBPPCS1WRDBUS_IN[117], PLBPPCS1WRDBUS[117]);
buf B_PLBPPCS1WRDBUS118 (PLBPPCS1WRDBUS_IN[118], PLBPPCS1WRDBUS[118]);
buf B_PLBPPCS1WRDBUS119 (PLBPPCS1WRDBUS_IN[119], PLBPPCS1WRDBUS[119]);
buf B_PLBPPCS1WRDBUS120 (PLBPPCS1WRDBUS_IN[120], PLBPPCS1WRDBUS[120]);
buf B_PLBPPCS1WRDBUS121 (PLBPPCS1WRDBUS_IN[121], PLBPPCS1WRDBUS[121]);
buf B_PLBPPCS1WRDBUS122 (PLBPPCS1WRDBUS_IN[122], PLBPPCS1WRDBUS[122]);
buf B_PLBPPCS1WRDBUS123 (PLBPPCS1WRDBUS_IN[123], PLBPPCS1WRDBUS[123]);
buf B_PLBPPCS1WRDBUS124 (PLBPPCS1WRDBUS_IN[124], PLBPPCS1WRDBUS[124]);
buf B_PLBPPCS1WRDBUS125 (PLBPPCS1WRDBUS_IN[125], PLBPPCS1WRDBUS[125]);
buf B_PLBPPCS1WRDBUS126 (PLBPPCS1WRDBUS_IN[126], PLBPPCS1WRDBUS[126]);
buf B_PLBPPCS1WRDBUS127 (PLBPPCS1WRDBUS_IN[127], PLBPPCS1WRDBUS[127]);
buf B_PLBPPCS1WRPENDPRI0 (PLBPPCS1WRPENDPRI_IN[0], PLBPPCS1WRPENDPRI[0]);
buf B_PLBPPCS1WRPENDPRI1 (PLBPPCS1WRPENDPRI_IN[1], PLBPPCS1WRPENDPRI[1]);
buf B_PLBPPCS1WRPENDREQ (PLBPPCS1WRPENDREQ_IN, PLBPPCS1WRPENDREQ);
buf B_PLBPPCS1WRPRIM (PLBPPCS1WRPRIM_IN, PLBPPCS1WRPRIM);
buf B_TIEDCRBASEADDR0 (TIEDCRBASEADDR_IN[0], TIEDCRBASEADDR[0]);
buf B_TIEDCRBASEADDR1 (TIEDCRBASEADDR_IN[1], TIEDCRBASEADDR[1]);
buf B_CPMC440CLK (CPMC440CLK_IN, CPMC440CLK);
buf B_CPMC440CLKEN (CPMC440CLKEN_IN, CPMC440CLKEN);
buf B_CPMC440CORECLOCKINACTIVE (CPMC440CORECLOCKINACTIVE_IN, CPMC440CORECLOCKINACTIVE);
buf B_CPMC440TIMERCLOCK (CPMC440TIMERCLOCK_IN, CPMC440TIMERCLOCK);
buf B_CPMFCMCLK (CPMFCMCLK_IN, CPMFCMCLK);
buf B_CPMINTERCONNECTCLK (CPMINTERCONNECTCLK_IN, CPMINTERCONNECTCLK);
buf B_CPMINTERCONNECTCLKEN (CPMINTERCONNECTCLKEN_IN, CPMINTERCONNECTCLKEN);
buf B_CPMMCCLK (CPMMCCLK_IN, CPMMCCLK);
buf B_DBGC440DEBUGHALT (DBGC440DEBUGHALT_IN, DBGC440DEBUGHALT);
buf B_DBGC440SYSTEMSTATUS0 (DBGC440SYSTEMSTATUS_IN[0], DBGC440SYSTEMSTATUS[0]);
buf B_DBGC440SYSTEMSTATUS1 (DBGC440SYSTEMSTATUS_IN[1], DBGC440SYSTEMSTATUS[1]);
buf B_DBGC440SYSTEMSTATUS2 (DBGC440SYSTEMSTATUS_IN[2], DBGC440SYSTEMSTATUS[2]);
buf B_DBGC440SYSTEMSTATUS3 (DBGC440SYSTEMSTATUS_IN[3], DBGC440SYSTEMSTATUS[3]);
buf B_DBGC440SYSTEMSTATUS4 (DBGC440SYSTEMSTATUS_IN[4], DBGC440SYSTEMSTATUS[4]);
buf B_DBGC440UNCONDDEBUGEVENT (DBGC440UNCONDDEBUGEVENT_IN, DBGC440UNCONDDEBUGEVENT);
buf B_DCRPPCDSABUS0 (DCRPPCDSABUS_IN[0], DCRPPCDSABUS[0]);
buf B_DCRPPCDSABUS1 (DCRPPCDSABUS_IN[1], DCRPPCDSABUS[1]);
buf B_DCRPPCDSABUS2 (DCRPPCDSABUS_IN[2], DCRPPCDSABUS[2]);
buf B_DCRPPCDSABUS3 (DCRPPCDSABUS_IN[3], DCRPPCDSABUS[3]);
buf B_DCRPPCDSABUS4 (DCRPPCDSABUS_IN[4], DCRPPCDSABUS[4]);
buf B_DCRPPCDSABUS5 (DCRPPCDSABUS_IN[5], DCRPPCDSABUS[5]);
buf B_DCRPPCDSABUS6 (DCRPPCDSABUS_IN[6], DCRPPCDSABUS[6]);
buf B_DCRPPCDSABUS7 (DCRPPCDSABUS_IN[7], DCRPPCDSABUS[7]);
buf B_DCRPPCDSABUS8 (DCRPPCDSABUS_IN[8], DCRPPCDSABUS[8]);
buf B_DCRPPCDSABUS9 (DCRPPCDSABUS_IN[9], DCRPPCDSABUS[9]);
buf B_DCRPPCDSDBUSOUT0 (DCRPPCDSDBUSOUT_IN[0], DCRPPCDSDBUSOUT[0]);
buf B_DCRPPCDSDBUSOUT1 (DCRPPCDSDBUSOUT_IN[1], DCRPPCDSDBUSOUT[1]);
buf B_DCRPPCDSDBUSOUT2 (DCRPPCDSDBUSOUT_IN[2], DCRPPCDSDBUSOUT[2]);
buf B_DCRPPCDSDBUSOUT3 (DCRPPCDSDBUSOUT_IN[3], DCRPPCDSDBUSOUT[3]);
buf B_DCRPPCDSDBUSOUT4 (DCRPPCDSDBUSOUT_IN[4], DCRPPCDSDBUSOUT[4]);
buf B_DCRPPCDSDBUSOUT5 (DCRPPCDSDBUSOUT_IN[5], DCRPPCDSDBUSOUT[5]);
buf B_DCRPPCDSDBUSOUT6 (DCRPPCDSDBUSOUT_IN[6], DCRPPCDSDBUSOUT[6]);
buf B_DCRPPCDSDBUSOUT7 (DCRPPCDSDBUSOUT_IN[7], DCRPPCDSDBUSOUT[7]);
buf B_DCRPPCDSDBUSOUT8 (DCRPPCDSDBUSOUT_IN[8], DCRPPCDSDBUSOUT[8]);
buf B_DCRPPCDSDBUSOUT9 (DCRPPCDSDBUSOUT_IN[9], DCRPPCDSDBUSOUT[9]);
buf B_DCRPPCDSDBUSOUT10 (DCRPPCDSDBUSOUT_IN[10], DCRPPCDSDBUSOUT[10]);
buf B_DCRPPCDSDBUSOUT11 (DCRPPCDSDBUSOUT_IN[11], DCRPPCDSDBUSOUT[11]);
buf B_DCRPPCDSDBUSOUT12 (DCRPPCDSDBUSOUT_IN[12], DCRPPCDSDBUSOUT[12]);
buf B_DCRPPCDSDBUSOUT13 (DCRPPCDSDBUSOUT_IN[13], DCRPPCDSDBUSOUT[13]);
buf B_DCRPPCDSDBUSOUT14 (DCRPPCDSDBUSOUT_IN[14], DCRPPCDSDBUSOUT[14]);
buf B_DCRPPCDSDBUSOUT15 (DCRPPCDSDBUSOUT_IN[15], DCRPPCDSDBUSOUT[15]);
buf B_DCRPPCDSDBUSOUT16 (DCRPPCDSDBUSOUT_IN[16], DCRPPCDSDBUSOUT[16]);
buf B_DCRPPCDSDBUSOUT17 (DCRPPCDSDBUSOUT_IN[17], DCRPPCDSDBUSOUT[17]);
buf B_DCRPPCDSDBUSOUT18 (DCRPPCDSDBUSOUT_IN[18], DCRPPCDSDBUSOUT[18]);
buf B_DCRPPCDSDBUSOUT19 (DCRPPCDSDBUSOUT_IN[19], DCRPPCDSDBUSOUT[19]);
buf B_DCRPPCDSDBUSOUT20 (DCRPPCDSDBUSOUT_IN[20], DCRPPCDSDBUSOUT[20]);
buf B_DCRPPCDSDBUSOUT21 (DCRPPCDSDBUSOUT_IN[21], DCRPPCDSDBUSOUT[21]);
buf B_DCRPPCDSDBUSOUT22 (DCRPPCDSDBUSOUT_IN[22], DCRPPCDSDBUSOUT[22]);
buf B_DCRPPCDSDBUSOUT23 (DCRPPCDSDBUSOUT_IN[23], DCRPPCDSDBUSOUT[23]);
buf B_DCRPPCDSDBUSOUT24 (DCRPPCDSDBUSOUT_IN[24], DCRPPCDSDBUSOUT[24]);
buf B_DCRPPCDSDBUSOUT25 (DCRPPCDSDBUSOUT_IN[25], DCRPPCDSDBUSOUT[25]);
buf B_DCRPPCDSDBUSOUT26 (DCRPPCDSDBUSOUT_IN[26], DCRPPCDSDBUSOUT[26]);
buf B_DCRPPCDSDBUSOUT27 (DCRPPCDSDBUSOUT_IN[27], DCRPPCDSDBUSOUT[27]);
buf B_DCRPPCDSDBUSOUT28 (DCRPPCDSDBUSOUT_IN[28], DCRPPCDSDBUSOUT[28]);
buf B_DCRPPCDSDBUSOUT29 (DCRPPCDSDBUSOUT_IN[29], DCRPPCDSDBUSOUT[29]);
buf B_DCRPPCDSDBUSOUT30 (DCRPPCDSDBUSOUT_IN[30], DCRPPCDSDBUSOUT[30]);
buf B_DCRPPCDSDBUSOUT31 (DCRPPCDSDBUSOUT_IN[31], DCRPPCDSDBUSOUT[31]);
buf B_DCRPPCDSREAD (DCRPPCDSREAD_IN, DCRPPCDSREAD);
buf B_DCRPPCDSWRITE (DCRPPCDSWRITE_IN, DCRPPCDSWRITE);
buf B_EICC440CRITIRQ (EICC440CRITIRQ_IN, EICC440CRITIRQ);
buf B_EICC440EXTIRQ (EICC440EXTIRQ_IN, EICC440EXTIRQ);
buf B_FCMAPUCONFIRMINSTR (FCMAPUCONFIRMINSTR_IN, FCMAPUCONFIRMINSTR);
buf B_FCMAPUCR0 (FCMAPUCR_IN[0], FCMAPUCR[0]);
buf B_FCMAPUCR1 (FCMAPUCR_IN[1], FCMAPUCR[1]);
buf B_FCMAPUCR2 (FCMAPUCR_IN[2], FCMAPUCR[2]);
buf B_FCMAPUCR3 (FCMAPUCR_IN[3], FCMAPUCR[3]);
buf B_FCMAPUDONE (FCMAPUDONE_IN, FCMAPUDONE);
buf B_FCMAPUEXCEPTION (FCMAPUEXCEPTION_IN, FCMAPUEXCEPTION);
buf B_FCMAPUFPSCRFEX (FCMAPUFPSCRFEX_IN, FCMAPUFPSCRFEX);
buf B_FCMAPURESULT0 (FCMAPURESULT_IN[0], FCMAPURESULT[0]);
buf B_FCMAPURESULT1 (FCMAPURESULT_IN[1], FCMAPURESULT[1]);
buf B_FCMAPURESULT2 (FCMAPURESULT_IN[2], FCMAPURESULT[2]);
buf B_FCMAPURESULT3 (FCMAPURESULT_IN[3], FCMAPURESULT[3]);
buf B_FCMAPURESULT4 (FCMAPURESULT_IN[4], FCMAPURESULT[4]);
buf B_FCMAPURESULT5 (FCMAPURESULT_IN[5], FCMAPURESULT[5]);
buf B_FCMAPURESULT6 (FCMAPURESULT_IN[6], FCMAPURESULT[6]);
buf B_FCMAPURESULT7 (FCMAPURESULT_IN[7], FCMAPURESULT[7]);
buf B_FCMAPURESULT8 (FCMAPURESULT_IN[8], FCMAPURESULT[8]);
buf B_FCMAPURESULT9 (FCMAPURESULT_IN[9], FCMAPURESULT[9]);
buf B_FCMAPURESULT10 (FCMAPURESULT_IN[10], FCMAPURESULT[10]);
buf B_FCMAPURESULT11 (FCMAPURESULT_IN[11], FCMAPURESULT[11]);
buf B_FCMAPURESULT12 (FCMAPURESULT_IN[12], FCMAPURESULT[12]);
buf B_FCMAPURESULT13 (FCMAPURESULT_IN[13], FCMAPURESULT[13]);
buf B_FCMAPURESULT14 (FCMAPURESULT_IN[14], FCMAPURESULT[14]);
buf B_FCMAPURESULT15 (FCMAPURESULT_IN[15], FCMAPURESULT[15]);
buf B_FCMAPURESULT16 (FCMAPURESULT_IN[16], FCMAPURESULT[16]);
buf B_FCMAPURESULT17 (FCMAPURESULT_IN[17], FCMAPURESULT[17]);
buf B_FCMAPURESULT18 (FCMAPURESULT_IN[18], FCMAPURESULT[18]);
buf B_FCMAPURESULT19 (FCMAPURESULT_IN[19], FCMAPURESULT[19]);
buf B_FCMAPURESULT20 (FCMAPURESULT_IN[20], FCMAPURESULT[20]);
buf B_FCMAPURESULT21 (FCMAPURESULT_IN[21], FCMAPURESULT[21]);
buf B_FCMAPURESULT22 (FCMAPURESULT_IN[22], FCMAPURESULT[22]);
buf B_FCMAPURESULT23 (FCMAPURESULT_IN[23], FCMAPURESULT[23]);
buf B_FCMAPURESULT24 (FCMAPURESULT_IN[24], FCMAPURESULT[24]);
buf B_FCMAPURESULT25 (FCMAPURESULT_IN[25], FCMAPURESULT[25]);
buf B_FCMAPURESULT26 (FCMAPURESULT_IN[26], FCMAPURESULT[26]);
buf B_FCMAPURESULT27 (FCMAPURESULT_IN[27], FCMAPURESULT[27]);
buf B_FCMAPURESULT28 (FCMAPURESULT_IN[28], FCMAPURESULT[28]);
buf B_FCMAPURESULT29 (FCMAPURESULT_IN[29], FCMAPURESULT[29]);
buf B_FCMAPURESULT30 (FCMAPURESULT_IN[30], FCMAPURESULT[30]);
buf B_FCMAPURESULT31 (FCMAPURESULT_IN[31], FCMAPURESULT[31]);
buf B_FCMAPURESULTVALID (FCMAPURESULTVALID_IN, FCMAPURESULTVALID);
buf B_FCMAPUSLEEPNOTREADY (FCMAPUSLEEPNOTREADY_IN, FCMAPUSLEEPNOTREADY);
buf B_FCMAPUSTOREDATA0 (FCMAPUSTOREDATA_IN[0], FCMAPUSTOREDATA[0]);
buf B_FCMAPUSTOREDATA1 (FCMAPUSTOREDATA_IN[1], FCMAPUSTOREDATA[1]);
buf B_FCMAPUSTOREDATA2 (FCMAPUSTOREDATA_IN[2], FCMAPUSTOREDATA[2]);
buf B_FCMAPUSTOREDATA3 (FCMAPUSTOREDATA_IN[3], FCMAPUSTOREDATA[3]);
buf B_FCMAPUSTOREDATA4 (FCMAPUSTOREDATA_IN[4], FCMAPUSTOREDATA[4]);
buf B_FCMAPUSTOREDATA5 (FCMAPUSTOREDATA_IN[5], FCMAPUSTOREDATA[5]);
buf B_FCMAPUSTOREDATA6 (FCMAPUSTOREDATA_IN[6], FCMAPUSTOREDATA[6]);
buf B_FCMAPUSTOREDATA7 (FCMAPUSTOREDATA_IN[7], FCMAPUSTOREDATA[7]);
buf B_FCMAPUSTOREDATA8 (FCMAPUSTOREDATA_IN[8], FCMAPUSTOREDATA[8]);
buf B_FCMAPUSTOREDATA9 (FCMAPUSTOREDATA_IN[9], FCMAPUSTOREDATA[9]);
buf B_FCMAPUSTOREDATA10 (FCMAPUSTOREDATA_IN[10], FCMAPUSTOREDATA[10]);
buf B_FCMAPUSTOREDATA11 (FCMAPUSTOREDATA_IN[11], FCMAPUSTOREDATA[11]);
buf B_FCMAPUSTOREDATA12 (FCMAPUSTOREDATA_IN[12], FCMAPUSTOREDATA[12]);
buf B_FCMAPUSTOREDATA13 (FCMAPUSTOREDATA_IN[13], FCMAPUSTOREDATA[13]);
buf B_FCMAPUSTOREDATA14 (FCMAPUSTOREDATA_IN[14], FCMAPUSTOREDATA[14]);
buf B_FCMAPUSTOREDATA15 (FCMAPUSTOREDATA_IN[15], FCMAPUSTOREDATA[15]);
buf B_FCMAPUSTOREDATA16 (FCMAPUSTOREDATA_IN[16], FCMAPUSTOREDATA[16]);
buf B_FCMAPUSTOREDATA17 (FCMAPUSTOREDATA_IN[17], FCMAPUSTOREDATA[17]);
buf B_FCMAPUSTOREDATA18 (FCMAPUSTOREDATA_IN[18], FCMAPUSTOREDATA[18]);
buf B_FCMAPUSTOREDATA19 (FCMAPUSTOREDATA_IN[19], FCMAPUSTOREDATA[19]);
buf B_FCMAPUSTOREDATA20 (FCMAPUSTOREDATA_IN[20], FCMAPUSTOREDATA[20]);
buf B_FCMAPUSTOREDATA21 (FCMAPUSTOREDATA_IN[21], FCMAPUSTOREDATA[21]);
buf B_FCMAPUSTOREDATA22 (FCMAPUSTOREDATA_IN[22], FCMAPUSTOREDATA[22]);
buf B_FCMAPUSTOREDATA23 (FCMAPUSTOREDATA_IN[23], FCMAPUSTOREDATA[23]);
buf B_FCMAPUSTOREDATA24 (FCMAPUSTOREDATA_IN[24], FCMAPUSTOREDATA[24]);
buf B_FCMAPUSTOREDATA25 (FCMAPUSTOREDATA_IN[25], FCMAPUSTOREDATA[25]);
buf B_FCMAPUSTOREDATA26 (FCMAPUSTOREDATA_IN[26], FCMAPUSTOREDATA[26]);
buf B_FCMAPUSTOREDATA27 (FCMAPUSTOREDATA_IN[27], FCMAPUSTOREDATA[27]);
buf B_FCMAPUSTOREDATA28 (FCMAPUSTOREDATA_IN[28], FCMAPUSTOREDATA[28]);
buf B_FCMAPUSTOREDATA29 (FCMAPUSTOREDATA_IN[29], FCMAPUSTOREDATA[29]);
buf B_FCMAPUSTOREDATA30 (FCMAPUSTOREDATA_IN[30], FCMAPUSTOREDATA[30]);
buf B_FCMAPUSTOREDATA31 (FCMAPUSTOREDATA_IN[31], FCMAPUSTOREDATA[31]);
buf B_FCMAPUSTOREDATA32 (FCMAPUSTOREDATA_IN[32], FCMAPUSTOREDATA[32]);
buf B_FCMAPUSTOREDATA33 (FCMAPUSTOREDATA_IN[33], FCMAPUSTOREDATA[33]);
buf B_FCMAPUSTOREDATA34 (FCMAPUSTOREDATA_IN[34], FCMAPUSTOREDATA[34]);
buf B_FCMAPUSTOREDATA35 (FCMAPUSTOREDATA_IN[35], FCMAPUSTOREDATA[35]);
buf B_FCMAPUSTOREDATA36 (FCMAPUSTOREDATA_IN[36], FCMAPUSTOREDATA[36]);
buf B_FCMAPUSTOREDATA37 (FCMAPUSTOREDATA_IN[37], FCMAPUSTOREDATA[37]);
buf B_FCMAPUSTOREDATA38 (FCMAPUSTOREDATA_IN[38], FCMAPUSTOREDATA[38]);
buf B_FCMAPUSTOREDATA39 (FCMAPUSTOREDATA_IN[39], FCMAPUSTOREDATA[39]);
buf B_FCMAPUSTOREDATA40 (FCMAPUSTOREDATA_IN[40], FCMAPUSTOREDATA[40]);
buf B_FCMAPUSTOREDATA41 (FCMAPUSTOREDATA_IN[41], FCMAPUSTOREDATA[41]);
buf B_FCMAPUSTOREDATA42 (FCMAPUSTOREDATA_IN[42], FCMAPUSTOREDATA[42]);
buf B_FCMAPUSTOREDATA43 (FCMAPUSTOREDATA_IN[43], FCMAPUSTOREDATA[43]);
buf B_FCMAPUSTOREDATA44 (FCMAPUSTOREDATA_IN[44], FCMAPUSTOREDATA[44]);
buf B_FCMAPUSTOREDATA45 (FCMAPUSTOREDATA_IN[45], FCMAPUSTOREDATA[45]);
buf B_FCMAPUSTOREDATA46 (FCMAPUSTOREDATA_IN[46], FCMAPUSTOREDATA[46]);
buf B_FCMAPUSTOREDATA47 (FCMAPUSTOREDATA_IN[47], FCMAPUSTOREDATA[47]);
buf B_FCMAPUSTOREDATA48 (FCMAPUSTOREDATA_IN[48], FCMAPUSTOREDATA[48]);
buf B_FCMAPUSTOREDATA49 (FCMAPUSTOREDATA_IN[49], FCMAPUSTOREDATA[49]);
buf B_FCMAPUSTOREDATA50 (FCMAPUSTOREDATA_IN[50], FCMAPUSTOREDATA[50]);
buf B_FCMAPUSTOREDATA51 (FCMAPUSTOREDATA_IN[51], FCMAPUSTOREDATA[51]);
buf B_FCMAPUSTOREDATA52 (FCMAPUSTOREDATA_IN[52], FCMAPUSTOREDATA[52]);
buf B_FCMAPUSTOREDATA53 (FCMAPUSTOREDATA_IN[53], FCMAPUSTOREDATA[53]);
buf B_FCMAPUSTOREDATA54 (FCMAPUSTOREDATA_IN[54], FCMAPUSTOREDATA[54]);
buf B_FCMAPUSTOREDATA55 (FCMAPUSTOREDATA_IN[55], FCMAPUSTOREDATA[55]);
buf B_FCMAPUSTOREDATA56 (FCMAPUSTOREDATA_IN[56], FCMAPUSTOREDATA[56]);
buf B_FCMAPUSTOREDATA57 (FCMAPUSTOREDATA_IN[57], FCMAPUSTOREDATA[57]);
buf B_FCMAPUSTOREDATA58 (FCMAPUSTOREDATA_IN[58], FCMAPUSTOREDATA[58]);
buf B_FCMAPUSTOREDATA59 (FCMAPUSTOREDATA_IN[59], FCMAPUSTOREDATA[59]);
buf B_FCMAPUSTOREDATA60 (FCMAPUSTOREDATA_IN[60], FCMAPUSTOREDATA[60]);
buf B_FCMAPUSTOREDATA61 (FCMAPUSTOREDATA_IN[61], FCMAPUSTOREDATA[61]);
buf B_FCMAPUSTOREDATA62 (FCMAPUSTOREDATA_IN[62], FCMAPUSTOREDATA[62]);
buf B_FCMAPUSTOREDATA63 (FCMAPUSTOREDATA_IN[63], FCMAPUSTOREDATA[63]);
buf B_FCMAPUSTOREDATA64 (FCMAPUSTOREDATA_IN[64], FCMAPUSTOREDATA[64]);
buf B_FCMAPUSTOREDATA65 (FCMAPUSTOREDATA_IN[65], FCMAPUSTOREDATA[65]);
buf B_FCMAPUSTOREDATA66 (FCMAPUSTOREDATA_IN[66], FCMAPUSTOREDATA[66]);
buf B_FCMAPUSTOREDATA67 (FCMAPUSTOREDATA_IN[67], FCMAPUSTOREDATA[67]);
buf B_FCMAPUSTOREDATA68 (FCMAPUSTOREDATA_IN[68], FCMAPUSTOREDATA[68]);
buf B_FCMAPUSTOREDATA69 (FCMAPUSTOREDATA_IN[69], FCMAPUSTOREDATA[69]);
buf B_FCMAPUSTOREDATA70 (FCMAPUSTOREDATA_IN[70], FCMAPUSTOREDATA[70]);
buf B_FCMAPUSTOREDATA71 (FCMAPUSTOREDATA_IN[71], FCMAPUSTOREDATA[71]);
buf B_FCMAPUSTOREDATA72 (FCMAPUSTOREDATA_IN[72], FCMAPUSTOREDATA[72]);
buf B_FCMAPUSTOREDATA73 (FCMAPUSTOREDATA_IN[73], FCMAPUSTOREDATA[73]);
buf B_FCMAPUSTOREDATA74 (FCMAPUSTOREDATA_IN[74], FCMAPUSTOREDATA[74]);
buf B_FCMAPUSTOREDATA75 (FCMAPUSTOREDATA_IN[75], FCMAPUSTOREDATA[75]);
buf B_FCMAPUSTOREDATA76 (FCMAPUSTOREDATA_IN[76], FCMAPUSTOREDATA[76]);
buf B_FCMAPUSTOREDATA77 (FCMAPUSTOREDATA_IN[77], FCMAPUSTOREDATA[77]);
buf B_FCMAPUSTOREDATA78 (FCMAPUSTOREDATA_IN[78], FCMAPUSTOREDATA[78]);
buf B_FCMAPUSTOREDATA79 (FCMAPUSTOREDATA_IN[79], FCMAPUSTOREDATA[79]);
buf B_FCMAPUSTOREDATA80 (FCMAPUSTOREDATA_IN[80], FCMAPUSTOREDATA[80]);
buf B_FCMAPUSTOREDATA81 (FCMAPUSTOREDATA_IN[81], FCMAPUSTOREDATA[81]);
buf B_FCMAPUSTOREDATA82 (FCMAPUSTOREDATA_IN[82], FCMAPUSTOREDATA[82]);
buf B_FCMAPUSTOREDATA83 (FCMAPUSTOREDATA_IN[83], FCMAPUSTOREDATA[83]);
buf B_FCMAPUSTOREDATA84 (FCMAPUSTOREDATA_IN[84], FCMAPUSTOREDATA[84]);
buf B_FCMAPUSTOREDATA85 (FCMAPUSTOREDATA_IN[85], FCMAPUSTOREDATA[85]);
buf B_FCMAPUSTOREDATA86 (FCMAPUSTOREDATA_IN[86], FCMAPUSTOREDATA[86]);
buf B_FCMAPUSTOREDATA87 (FCMAPUSTOREDATA_IN[87], FCMAPUSTOREDATA[87]);
buf B_FCMAPUSTOREDATA88 (FCMAPUSTOREDATA_IN[88], FCMAPUSTOREDATA[88]);
buf B_FCMAPUSTOREDATA89 (FCMAPUSTOREDATA_IN[89], FCMAPUSTOREDATA[89]);
buf B_FCMAPUSTOREDATA90 (FCMAPUSTOREDATA_IN[90], FCMAPUSTOREDATA[90]);
buf B_FCMAPUSTOREDATA91 (FCMAPUSTOREDATA_IN[91], FCMAPUSTOREDATA[91]);
buf B_FCMAPUSTOREDATA92 (FCMAPUSTOREDATA_IN[92], FCMAPUSTOREDATA[92]);
buf B_FCMAPUSTOREDATA93 (FCMAPUSTOREDATA_IN[93], FCMAPUSTOREDATA[93]);
buf B_FCMAPUSTOREDATA94 (FCMAPUSTOREDATA_IN[94], FCMAPUSTOREDATA[94]);
buf B_FCMAPUSTOREDATA95 (FCMAPUSTOREDATA_IN[95], FCMAPUSTOREDATA[95]);
buf B_FCMAPUSTOREDATA96 (FCMAPUSTOREDATA_IN[96], FCMAPUSTOREDATA[96]);
buf B_FCMAPUSTOREDATA97 (FCMAPUSTOREDATA_IN[97], FCMAPUSTOREDATA[97]);
buf B_FCMAPUSTOREDATA98 (FCMAPUSTOREDATA_IN[98], FCMAPUSTOREDATA[98]);
buf B_FCMAPUSTOREDATA99 (FCMAPUSTOREDATA_IN[99], FCMAPUSTOREDATA[99]);
buf B_FCMAPUSTOREDATA100 (FCMAPUSTOREDATA_IN[100], FCMAPUSTOREDATA[100]);
buf B_FCMAPUSTOREDATA101 (FCMAPUSTOREDATA_IN[101], FCMAPUSTOREDATA[101]);
buf B_FCMAPUSTOREDATA102 (FCMAPUSTOREDATA_IN[102], FCMAPUSTOREDATA[102]);
buf B_FCMAPUSTOREDATA103 (FCMAPUSTOREDATA_IN[103], FCMAPUSTOREDATA[103]);
buf B_FCMAPUSTOREDATA104 (FCMAPUSTOREDATA_IN[104], FCMAPUSTOREDATA[104]);
buf B_FCMAPUSTOREDATA105 (FCMAPUSTOREDATA_IN[105], FCMAPUSTOREDATA[105]);
buf B_FCMAPUSTOREDATA106 (FCMAPUSTOREDATA_IN[106], FCMAPUSTOREDATA[106]);
buf B_FCMAPUSTOREDATA107 (FCMAPUSTOREDATA_IN[107], FCMAPUSTOREDATA[107]);
buf B_FCMAPUSTOREDATA108 (FCMAPUSTOREDATA_IN[108], FCMAPUSTOREDATA[108]);
buf B_FCMAPUSTOREDATA109 (FCMAPUSTOREDATA_IN[109], FCMAPUSTOREDATA[109]);
buf B_FCMAPUSTOREDATA110 (FCMAPUSTOREDATA_IN[110], FCMAPUSTOREDATA[110]);
buf B_FCMAPUSTOREDATA111 (FCMAPUSTOREDATA_IN[111], FCMAPUSTOREDATA[111]);
buf B_FCMAPUSTOREDATA112 (FCMAPUSTOREDATA_IN[112], FCMAPUSTOREDATA[112]);
buf B_FCMAPUSTOREDATA113 (FCMAPUSTOREDATA_IN[113], FCMAPUSTOREDATA[113]);
buf B_FCMAPUSTOREDATA114 (FCMAPUSTOREDATA_IN[114], FCMAPUSTOREDATA[114]);
buf B_FCMAPUSTOREDATA115 (FCMAPUSTOREDATA_IN[115], FCMAPUSTOREDATA[115]);
buf B_FCMAPUSTOREDATA116 (FCMAPUSTOREDATA_IN[116], FCMAPUSTOREDATA[116]);
buf B_FCMAPUSTOREDATA117 (FCMAPUSTOREDATA_IN[117], FCMAPUSTOREDATA[117]);
buf B_FCMAPUSTOREDATA118 (FCMAPUSTOREDATA_IN[118], FCMAPUSTOREDATA[118]);
buf B_FCMAPUSTOREDATA119 (FCMAPUSTOREDATA_IN[119], FCMAPUSTOREDATA[119]);
buf B_FCMAPUSTOREDATA120 (FCMAPUSTOREDATA_IN[120], FCMAPUSTOREDATA[120]);
buf B_FCMAPUSTOREDATA121 (FCMAPUSTOREDATA_IN[121], FCMAPUSTOREDATA[121]);
buf B_FCMAPUSTOREDATA122 (FCMAPUSTOREDATA_IN[122], FCMAPUSTOREDATA[122]);
buf B_FCMAPUSTOREDATA123 (FCMAPUSTOREDATA_IN[123], FCMAPUSTOREDATA[123]);
buf B_FCMAPUSTOREDATA124 (FCMAPUSTOREDATA_IN[124], FCMAPUSTOREDATA[124]);
buf B_FCMAPUSTOREDATA125 (FCMAPUSTOREDATA_IN[125], FCMAPUSTOREDATA[125]);
buf B_FCMAPUSTOREDATA126 (FCMAPUSTOREDATA_IN[126], FCMAPUSTOREDATA[126]);
buf B_FCMAPUSTOREDATA127 (FCMAPUSTOREDATA_IN[127], FCMAPUSTOREDATA[127]);
buf B_JTGC440TCK (JTGC440TCK_IN, JTGC440TCK);
buf B_JTGC440TDI (JTGC440TDI_IN, JTGC440TDI);
buf B_JTGC440TMS (JTGC440TMS_IN, JTGC440TMS);
buf B_JTGC440TRSTNEG (JTGC440TRSTNEG_IN, JTGC440TRSTNEG);
buf B_MCMIADDRREADYTOACCEPT (MCMIADDRREADYTOACCEPT_IN, MCMIADDRREADYTOACCEPT);
buf B_MCMIREADDATA0 (MCMIREADDATA_IN[0], MCMIREADDATA[0]);
buf B_MCMIREADDATA1 (MCMIREADDATA_IN[1], MCMIREADDATA[1]);
buf B_MCMIREADDATA2 (MCMIREADDATA_IN[2], MCMIREADDATA[2]);
buf B_MCMIREADDATA3 (MCMIREADDATA_IN[3], MCMIREADDATA[3]);
buf B_MCMIREADDATA4 (MCMIREADDATA_IN[4], MCMIREADDATA[4]);
buf B_MCMIREADDATA5 (MCMIREADDATA_IN[5], MCMIREADDATA[5]);
buf B_MCMIREADDATA6 (MCMIREADDATA_IN[6], MCMIREADDATA[6]);
buf B_MCMIREADDATA7 (MCMIREADDATA_IN[7], MCMIREADDATA[7]);
buf B_MCMIREADDATA8 (MCMIREADDATA_IN[8], MCMIREADDATA[8]);
buf B_MCMIREADDATA9 (MCMIREADDATA_IN[9], MCMIREADDATA[9]);
buf B_MCMIREADDATA10 (MCMIREADDATA_IN[10], MCMIREADDATA[10]);
buf B_MCMIREADDATA11 (MCMIREADDATA_IN[11], MCMIREADDATA[11]);
buf B_MCMIREADDATA12 (MCMIREADDATA_IN[12], MCMIREADDATA[12]);
buf B_MCMIREADDATA13 (MCMIREADDATA_IN[13], MCMIREADDATA[13]);
buf B_MCMIREADDATA14 (MCMIREADDATA_IN[14], MCMIREADDATA[14]);
buf B_MCMIREADDATA15 (MCMIREADDATA_IN[15], MCMIREADDATA[15]);
buf B_MCMIREADDATA16 (MCMIREADDATA_IN[16], MCMIREADDATA[16]);
buf B_MCMIREADDATA17 (MCMIREADDATA_IN[17], MCMIREADDATA[17]);
buf B_MCMIREADDATA18 (MCMIREADDATA_IN[18], MCMIREADDATA[18]);
buf B_MCMIREADDATA19 (MCMIREADDATA_IN[19], MCMIREADDATA[19]);
buf B_MCMIREADDATA20 (MCMIREADDATA_IN[20], MCMIREADDATA[20]);
buf B_MCMIREADDATA21 (MCMIREADDATA_IN[21], MCMIREADDATA[21]);
buf B_MCMIREADDATA22 (MCMIREADDATA_IN[22], MCMIREADDATA[22]);
buf B_MCMIREADDATA23 (MCMIREADDATA_IN[23], MCMIREADDATA[23]);
buf B_MCMIREADDATA24 (MCMIREADDATA_IN[24], MCMIREADDATA[24]);
buf B_MCMIREADDATA25 (MCMIREADDATA_IN[25], MCMIREADDATA[25]);
buf B_MCMIREADDATA26 (MCMIREADDATA_IN[26], MCMIREADDATA[26]);
buf B_MCMIREADDATA27 (MCMIREADDATA_IN[27], MCMIREADDATA[27]);
buf B_MCMIREADDATA28 (MCMIREADDATA_IN[28], MCMIREADDATA[28]);
buf B_MCMIREADDATA29 (MCMIREADDATA_IN[29], MCMIREADDATA[29]);
buf B_MCMIREADDATA30 (MCMIREADDATA_IN[30], MCMIREADDATA[30]);
buf B_MCMIREADDATA31 (MCMIREADDATA_IN[31], MCMIREADDATA[31]);
buf B_MCMIREADDATA32 (MCMIREADDATA_IN[32], MCMIREADDATA[32]);
buf B_MCMIREADDATA33 (MCMIREADDATA_IN[33], MCMIREADDATA[33]);
buf B_MCMIREADDATA34 (MCMIREADDATA_IN[34], MCMIREADDATA[34]);
buf B_MCMIREADDATA35 (MCMIREADDATA_IN[35], MCMIREADDATA[35]);
buf B_MCMIREADDATA36 (MCMIREADDATA_IN[36], MCMIREADDATA[36]);
buf B_MCMIREADDATA37 (MCMIREADDATA_IN[37], MCMIREADDATA[37]);
buf B_MCMIREADDATA38 (MCMIREADDATA_IN[38], MCMIREADDATA[38]);
buf B_MCMIREADDATA39 (MCMIREADDATA_IN[39], MCMIREADDATA[39]);
buf B_MCMIREADDATA40 (MCMIREADDATA_IN[40], MCMIREADDATA[40]);
buf B_MCMIREADDATA41 (MCMIREADDATA_IN[41], MCMIREADDATA[41]);
buf B_MCMIREADDATA42 (MCMIREADDATA_IN[42], MCMIREADDATA[42]);
buf B_MCMIREADDATA43 (MCMIREADDATA_IN[43], MCMIREADDATA[43]);
buf B_MCMIREADDATA44 (MCMIREADDATA_IN[44], MCMIREADDATA[44]);
buf B_MCMIREADDATA45 (MCMIREADDATA_IN[45], MCMIREADDATA[45]);
buf B_MCMIREADDATA46 (MCMIREADDATA_IN[46], MCMIREADDATA[46]);
buf B_MCMIREADDATA47 (MCMIREADDATA_IN[47], MCMIREADDATA[47]);
buf B_MCMIREADDATA48 (MCMIREADDATA_IN[48], MCMIREADDATA[48]);
buf B_MCMIREADDATA49 (MCMIREADDATA_IN[49], MCMIREADDATA[49]);
buf B_MCMIREADDATA50 (MCMIREADDATA_IN[50], MCMIREADDATA[50]);
buf B_MCMIREADDATA51 (MCMIREADDATA_IN[51], MCMIREADDATA[51]);
buf B_MCMIREADDATA52 (MCMIREADDATA_IN[52], MCMIREADDATA[52]);
buf B_MCMIREADDATA53 (MCMIREADDATA_IN[53], MCMIREADDATA[53]);
buf B_MCMIREADDATA54 (MCMIREADDATA_IN[54], MCMIREADDATA[54]);
buf B_MCMIREADDATA55 (MCMIREADDATA_IN[55], MCMIREADDATA[55]);
buf B_MCMIREADDATA56 (MCMIREADDATA_IN[56], MCMIREADDATA[56]);
buf B_MCMIREADDATA57 (MCMIREADDATA_IN[57], MCMIREADDATA[57]);
buf B_MCMIREADDATA58 (MCMIREADDATA_IN[58], MCMIREADDATA[58]);
buf B_MCMIREADDATA59 (MCMIREADDATA_IN[59], MCMIREADDATA[59]);
buf B_MCMIREADDATA60 (MCMIREADDATA_IN[60], MCMIREADDATA[60]);
buf B_MCMIREADDATA61 (MCMIREADDATA_IN[61], MCMIREADDATA[61]);
buf B_MCMIREADDATA62 (MCMIREADDATA_IN[62], MCMIREADDATA[62]);
buf B_MCMIREADDATA63 (MCMIREADDATA_IN[63], MCMIREADDATA[63]);
buf B_MCMIREADDATA64 (MCMIREADDATA_IN[64], MCMIREADDATA[64]);
buf B_MCMIREADDATA65 (MCMIREADDATA_IN[65], MCMIREADDATA[65]);
buf B_MCMIREADDATA66 (MCMIREADDATA_IN[66], MCMIREADDATA[66]);
buf B_MCMIREADDATA67 (MCMIREADDATA_IN[67], MCMIREADDATA[67]);
buf B_MCMIREADDATA68 (MCMIREADDATA_IN[68], MCMIREADDATA[68]);
buf B_MCMIREADDATA69 (MCMIREADDATA_IN[69], MCMIREADDATA[69]);
buf B_MCMIREADDATA70 (MCMIREADDATA_IN[70], MCMIREADDATA[70]);
buf B_MCMIREADDATA71 (MCMIREADDATA_IN[71], MCMIREADDATA[71]);
buf B_MCMIREADDATA72 (MCMIREADDATA_IN[72], MCMIREADDATA[72]);
buf B_MCMIREADDATA73 (MCMIREADDATA_IN[73], MCMIREADDATA[73]);
buf B_MCMIREADDATA74 (MCMIREADDATA_IN[74], MCMIREADDATA[74]);
buf B_MCMIREADDATA75 (MCMIREADDATA_IN[75], MCMIREADDATA[75]);
buf B_MCMIREADDATA76 (MCMIREADDATA_IN[76], MCMIREADDATA[76]);
buf B_MCMIREADDATA77 (MCMIREADDATA_IN[77], MCMIREADDATA[77]);
buf B_MCMIREADDATA78 (MCMIREADDATA_IN[78], MCMIREADDATA[78]);
buf B_MCMIREADDATA79 (MCMIREADDATA_IN[79], MCMIREADDATA[79]);
buf B_MCMIREADDATA80 (MCMIREADDATA_IN[80], MCMIREADDATA[80]);
buf B_MCMIREADDATA81 (MCMIREADDATA_IN[81], MCMIREADDATA[81]);
buf B_MCMIREADDATA82 (MCMIREADDATA_IN[82], MCMIREADDATA[82]);
buf B_MCMIREADDATA83 (MCMIREADDATA_IN[83], MCMIREADDATA[83]);
buf B_MCMIREADDATA84 (MCMIREADDATA_IN[84], MCMIREADDATA[84]);
buf B_MCMIREADDATA85 (MCMIREADDATA_IN[85], MCMIREADDATA[85]);
buf B_MCMIREADDATA86 (MCMIREADDATA_IN[86], MCMIREADDATA[86]);
buf B_MCMIREADDATA87 (MCMIREADDATA_IN[87], MCMIREADDATA[87]);
buf B_MCMIREADDATA88 (MCMIREADDATA_IN[88], MCMIREADDATA[88]);
buf B_MCMIREADDATA89 (MCMIREADDATA_IN[89], MCMIREADDATA[89]);
buf B_MCMIREADDATA90 (MCMIREADDATA_IN[90], MCMIREADDATA[90]);
buf B_MCMIREADDATA91 (MCMIREADDATA_IN[91], MCMIREADDATA[91]);
buf B_MCMIREADDATA92 (MCMIREADDATA_IN[92], MCMIREADDATA[92]);
buf B_MCMIREADDATA93 (MCMIREADDATA_IN[93], MCMIREADDATA[93]);
buf B_MCMIREADDATA94 (MCMIREADDATA_IN[94], MCMIREADDATA[94]);
buf B_MCMIREADDATA95 (MCMIREADDATA_IN[95], MCMIREADDATA[95]);
buf B_MCMIREADDATA96 (MCMIREADDATA_IN[96], MCMIREADDATA[96]);
buf B_MCMIREADDATA97 (MCMIREADDATA_IN[97], MCMIREADDATA[97]);
buf B_MCMIREADDATA98 (MCMIREADDATA_IN[98], MCMIREADDATA[98]);
buf B_MCMIREADDATA99 (MCMIREADDATA_IN[99], MCMIREADDATA[99]);
buf B_MCMIREADDATA100 (MCMIREADDATA_IN[100], MCMIREADDATA[100]);
buf B_MCMIREADDATA101 (MCMIREADDATA_IN[101], MCMIREADDATA[101]);
buf B_MCMIREADDATA102 (MCMIREADDATA_IN[102], MCMIREADDATA[102]);
buf B_MCMIREADDATA103 (MCMIREADDATA_IN[103], MCMIREADDATA[103]);
buf B_MCMIREADDATA104 (MCMIREADDATA_IN[104], MCMIREADDATA[104]);
buf B_MCMIREADDATA105 (MCMIREADDATA_IN[105], MCMIREADDATA[105]);
buf B_MCMIREADDATA106 (MCMIREADDATA_IN[106], MCMIREADDATA[106]);
buf B_MCMIREADDATA107 (MCMIREADDATA_IN[107], MCMIREADDATA[107]);
buf B_MCMIREADDATA108 (MCMIREADDATA_IN[108], MCMIREADDATA[108]);
buf B_MCMIREADDATA109 (MCMIREADDATA_IN[109], MCMIREADDATA[109]);
buf B_MCMIREADDATA110 (MCMIREADDATA_IN[110], MCMIREADDATA[110]);
buf B_MCMIREADDATA111 (MCMIREADDATA_IN[111], MCMIREADDATA[111]);
buf B_MCMIREADDATA112 (MCMIREADDATA_IN[112], MCMIREADDATA[112]);
buf B_MCMIREADDATA113 (MCMIREADDATA_IN[113], MCMIREADDATA[113]);
buf B_MCMIREADDATA114 (MCMIREADDATA_IN[114], MCMIREADDATA[114]);
buf B_MCMIREADDATA115 (MCMIREADDATA_IN[115], MCMIREADDATA[115]);
buf B_MCMIREADDATA116 (MCMIREADDATA_IN[116], MCMIREADDATA[116]);
buf B_MCMIREADDATA117 (MCMIREADDATA_IN[117], MCMIREADDATA[117]);
buf B_MCMIREADDATA118 (MCMIREADDATA_IN[118], MCMIREADDATA[118]);
buf B_MCMIREADDATA119 (MCMIREADDATA_IN[119], MCMIREADDATA[119]);
buf B_MCMIREADDATA120 (MCMIREADDATA_IN[120], MCMIREADDATA[120]);
buf B_MCMIREADDATA121 (MCMIREADDATA_IN[121], MCMIREADDATA[121]);
buf B_MCMIREADDATA122 (MCMIREADDATA_IN[122], MCMIREADDATA[122]);
buf B_MCMIREADDATA123 (MCMIREADDATA_IN[123], MCMIREADDATA[123]);
buf B_MCMIREADDATA124 (MCMIREADDATA_IN[124], MCMIREADDATA[124]);
buf B_MCMIREADDATA125 (MCMIREADDATA_IN[125], MCMIREADDATA[125]);
buf B_MCMIREADDATA126 (MCMIREADDATA_IN[126], MCMIREADDATA[126]);
buf B_MCMIREADDATA127 (MCMIREADDATA_IN[127], MCMIREADDATA[127]);
buf B_MCMIREADDATAERR (MCMIREADDATAERR_IN, MCMIREADDATAERR);
buf B_MCMIREADDATAVALID (MCMIREADDATAVALID_IN, MCMIREADDATAVALID);
buf B_RSTC440RESETCHIP (RSTC440RESETCHIP_IN, RSTC440RESETCHIP);
buf B_RSTC440RESETCORE (RSTC440RESETCORE_IN, RSTC440RESETCORE);
buf B_RSTC440RESETSYSTEM (RSTC440RESETSYSTEM_IN, RSTC440RESETSYSTEM);
buf B_TIEC440DCURDLDCACHEPLBPRIO0 (TIEC440DCURDLDCACHEPLBPRIO_IN[0], TIEC440DCURDLDCACHEPLBPRIO[0]);
buf B_TIEC440DCURDLDCACHEPLBPRIO1 (TIEC440DCURDLDCACHEPLBPRIO_IN[1], TIEC440DCURDLDCACHEPLBPRIO[1]);
buf B_TIEC440DCURDNONCACHEPLBPRIO0 (TIEC440DCURDNONCACHEPLBPRIO_IN[0], TIEC440DCURDNONCACHEPLBPRIO[0]);
buf B_TIEC440DCURDNONCACHEPLBPRIO1 (TIEC440DCURDNONCACHEPLBPRIO_IN[1], TIEC440DCURDNONCACHEPLBPRIO[1]);
buf B_TIEC440DCURDTOUCHPLBPRIO0 (TIEC440DCURDTOUCHPLBPRIO_IN[0], TIEC440DCURDTOUCHPLBPRIO[0]);
buf B_TIEC440DCURDTOUCHPLBPRIO1 (TIEC440DCURDTOUCHPLBPRIO_IN[1], TIEC440DCURDTOUCHPLBPRIO[1]);
buf B_TIEC440DCURDURGENTPLBPRIO0 (TIEC440DCURDURGENTPLBPRIO_IN[0], TIEC440DCURDURGENTPLBPRIO[0]);
buf B_TIEC440DCURDURGENTPLBPRIO1 (TIEC440DCURDURGENTPLBPRIO_IN[1], TIEC440DCURDURGENTPLBPRIO[1]);
buf B_TIEC440DCUWRFLUSHPLBPRIO0 (TIEC440DCUWRFLUSHPLBPRIO_IN[0], TIEC440DCUWRFLUSHPLBPRIO[0]);
buf B_TIEC440DCUWRFLUSHPLBPRIO1 (TIEC440DCUWRFLUSHPLBPRIO_IN[1], TIEC440DCUWRFLUSHPLBPRIO[1]);
buf B_TIEC440DCUWRSTOREPLBPRIO0 (TIEC440DCUWRSTOREPLBPRIO_IN[0], TIEC440DCUWRSTOREPLBPRIO[0]);
buf B_TIEC440DCUWRSTOREPLBPRIO1 (TIEC440DCUWRSTOREPLBPRIO_IN[1], TIEC440DCUWRSTOREPLBPRIO[1]);
buf B_TIEC440DCUWRURGENTPLBPRIO0 (TIEC440DCUWRURGENTPLBPRIO_IN[0], TIEC440DCUWRURGENTPLBPRIO[0]);
buf B_TIEC440DCUWRURGENTPLBPRIO1 (TIEC440DCUWRURGENTPLBPRIO_IN[1], TIEC440DCUWRURGENTPLBPRIO[1]);
buf B_TIEC440ENDIANRESET (TIEC440ENDIANRESET_IN, TIEC440ENDIANRESET);
buf B_TIEC440ERPNRESET0 (TIEC440ERPNRESET_IN[0], TIEC440ERPNRESET[0]);
buf B_TIEC440ERPNRESET1 (TIEC440ERPNRESET_IN[1], TIEC440ERPNRESET[1]);
buf B_TIEC440ERPNRESET2 (TIEC440ERPNRESET_IN[2], TIEC440ERPNRESET[2]);
buf B_TIEC440ERPNRESET3 (TIEC440ERPNRESET_IN[3], TIEC440ERPNRESET[3]);
buf B_TIEC440ICURDFETCHPLBPRIO0 (TIEC440ICURDFETCHPLBPRIO_IN[0], TIEC440ICURDFETCHPLBPRIO[0]);
buf B_TIEC440ICURDFETCHPLBPRIO1 (TIEC440ICURDFETCHPLBPRIO_IN[1], TIEC440ICURDFETCHPLBPRIO[1]);
buf B_TIEC440ICURDSPECPLBPRIO0 (TIEC440ICURDSPECPLBPRIO_IN[0], TIEC440ICURDSPECPLBPRIO[0]);
buf B_TIEC440ICURDSPECPLBPRIO1 (TIEC440ICURDSPECPLBPRIO_IN[1], TIEC440ICURDSPECPLBPRIO[1]);
buf B_TIEC440ICURDTOUCHPLBPRIO0 (TIEC440ICURDTOUCHPLBPRIO_IN[0], TIEC440ICURDTOUCHPLBPRIO[0]);
buf B_TIEC440ICURDTOUCHPLBPRIO1 (TIEC440ICURDTOUCHPLBPRIO_IN[1], TIEC440ICURDTOUCHPLBPRIO[1]);
buf B_TIEC440PIR28 (TIEC440PIR_IN[28], TIEC440PIR[28]);
buf B_TIEC440PIR29 (TIEC440PIR_IN[29], TIEC440PIR[29]);
buf B_TIEC440PIR30 (TIEC440PIR_IN[30], TIEC440PIR[30]);
buf B_TIEC440PIR31 (TIEC440PIR_IN[31], TIEC440PIR[31]);
buf B_TIEC440PVR28 (TIEC440PVR_IN[28], TIEC440PVR[28]);
buf B_TIEC440PVR29 (TIEC440PVR_IN[29], TIEC440PVR[29]);
buf B_TIEC440PVR30 (TIEC440PVR_IN[30], TIEC440PVR[30]);
buf B_TIEC440PVR31 (TIEC440PVR_IN[31], TIEC440PVR[31]);
buf B_TIEC440USERRESET0 (TIEC440USERRESET_IN[0], TIEC440USERRESET[0]);
buf B_TIEC440USERRESET1 (TIEC440USERRESET_IN[1], TIEC440USERRESET[1]);
buf B_TIEC440USERRESET2 (TIEC440USERRESET_IN[2], TIEC440USERRESET[2]);
buf B_TIEC440USERRESET3 (TIEC440USERRESET_IN[3], TIEC440USERRESET[3]);
buf B_TRCC440TRACEDISABLE (TRCC440TRACEDISABLE_IN, TRCC440TRACEDISABLE);
buf B_TRCC440TRIGGEREVENTIN (TRCC440TRIGGEREVENTIN_IN, TRCC440TRIGGEREVENTIN);

wire APUFCMDECFPUOP_delay;
wire APUFCMDECLOAD_delay;
wire APUFCMDECNONAUTON_delay;
wire APUFCMDECSTORE_delay;
wire APUFCMDECUDIVALID_delay;
wire APUFCMENDIAN_delay;
wire APUFCMFLUSH_delay;
wire APUFCMINSTRVALID_delay;
wire APUFCMLOADDVALID_delay;
wire APUFCMMSRFE0_delay;
wire APUFCMMSRFE1_delay;
wire APUFCMNEXTINSTRREADY_delay;
wire APUFCMOPERANDVALID_delay;
wire APUFCMWRITEBACKOK_delay;
wire C440CPMCORESLEEPREQ_delay;
wire C440CPMDECIRPTREQ_delay;
wire C440CPMFITIRPTREQ_delay;
wire C440CPMMSRCE_delay;
wire C440CPMMSREE_delay;
wire C440CPMTIMERRESETREQ_delay;
wire C440CPMWDIRPTREQ_delay;
wire C440JTGTDOEN_delay;
wire C440JTGTDO_delay;
wire C440MACHINECHECK_delay;
wire C440RSTCHIPRESETREQ_delay;
wire C440RSTCORERESETREQ_delay;
wire C440RSTSYSTEMRESETREQ_delay;
wire C440TRCCYCLE_delay;
wire C440TRCTRIGGEREVENTOUT_delay;
wire DMA0LLRSTENGINEACK_delay;
wire DMA0LLRXDSTRDYN_delay;
wire DMA0LLTXEOFN_delay;
wire DMA0LLTXEOPN_delay;
wire DMA0LLTXSOFN_delay;
wire DMA0LLTXSOPN_delay;
wire DMA0LLTXSRCRDYN_delay;
wire DMA0RXIRQ_delay;
wire DMA0TXIRQ_delay;
wire DMA1LLRSTENGINEACK_delay;
wire DMA1LLRXDSTRDYN_delay;
wire DMA1LLTXEOFN_delay;
wire DMA1LLTXEOPN_delay;
wire DMA1LLTXSOFN_delay;
wire DMA1LLTXSOPN_delay;
wire DMA1LLTXSRCRDYN_delay;
wire DMA1RXIRQ_delay;
wire DMA1TXIRQ_delay;
wire DMA2LLRSTENGINEACK_delay;
wire DMA2LLRXDSTRDYN_delay;
wire DMA2LLTXEOFN_delay;
wire DMA2LLTXEOPN_delay;
wire DMA2LLTXSOFN_delay;
wire DMA2LLTXSOPN_delay;
wire DMA2LLTXSRCRDYN_delay;
wire DMA2RXIRQ_delay;
wire DMA2TXIRQ_delay;
wire DMA3LLRSTENGINEACK_delay;
wire DMA3LLRXDSTRDYN_delay;
wire DMA3LLTXEOFN_delay;
wire DMA3LLTXEOPN_delay;
wire DMA3LLTXSOFN_delay;
wire DMA3LLTXSOPN_delay;
wire DMA3LLTXSRCRDYN_delay;
wire DMA3RXIRQ_delay;
wire DMA3TXIRQ_delay;
wire MIMCADDRESSVALID_delay;
wire MIMCBANKCONFLICT_delay;
wire MIMCREADNOTWRITE_delay;
wire MIMCROWCONFLICT_delay;
wire MIMCWRITEDATAVALID_delay;
wire PPCCPMINTERCONNECTBUSY_delay;
wire PPCDMDCRREAD_delay;
wire PPCDMDCRWRITE_delay;
wire PPCDSDCRACK_delay;
wire PPCDSDCRTIMEOUTWAIT_delay;
wire PPCEICINTERCONNECTIRQ_delay;
wire PPCMPLBABORT_delay;
wire PPCMPLBBUSLOCK_delay;
wire PPCMPLBLOCKERR_delay;
wire PPCMPLBRDBURST_delay;
wire PPCMPLBREQUEST_delay;
wire PPCMPLBRNW_delay;
wire PPCMPLBWRBURST_delay;
wire PPCS0PLBADDRACK_delay;
wire PPCS0PLBRDBTERM_delay;
wire PPCS0PLBRDCOMP_delay;
wire PPCS0PLBRDDACK_delay;
wire PPCS0PLBREARBITRATE_delay;
wire PPCS0PLBWAIT_delay;
wire PPCS0PLBWRBTERM_delay;
wire PPCS0PLBWRCOMP_delay;
wire PPCS0PLBWRDACK_delay;
wire PPCS1PLBADDRACK_delay;
wire PPCS1PLBRDBTERM_delay;
wire PPCS1PLBRDCOMP_delay;
wire PPCS1PLBRDDACK_delay;
wire PPCS1PLBREARBITRATE_delay;
wire PPCS1PLBWAIT_delay;
wire PPCS1PLBWRBTERM_delay;
wire PPCS1PLBWRCOMP_delay;
wire PPCS1PLBWRDACK_delay;
wire [0:127] APUFCMLOADDATA_delay;
wire [0:127] MIMCWRITEDATA_delay;
wire [0:127] PPCMPLBWRDBUS_delay;
wire [0:127] PPCS0PLBRDDBUS_delay;
wire [0:127] PPCS1PLBRDDBUS_delay;
wire [0:13] C440TRCTRIGGEREVENTTYPE_delay;
wire [0:15] MIMCBYTEENABLE_delay;
wire [0:15] PPCMPLBBE_delay;
wire [0:15] PPCMPLBTATTRIBUTE_delay;
wire [0:1] PPCMPLBPRIORITY_delay;
wire [0:1] PPCS0PLBSSIZE_delay;
wire [0:1] PPCS1PLBSSIZE_delay;
wire [0:2] APUFCMDECLDSTXFERSIZE_delay;
wire [0:2] C440TRCBRANCHSTATUS_delay;
wire [0:2] PPCMPLBTYPE_delay;
wire [0:31] APUFCMINSTRUCTION_delay;
wire [0:31] APUFCMRADATA_delay;
wire [0:31] APUFCMRBDATA_delay;
wire [0:31] DMA0LLTXD_delay;
wire [0:31] DMA1LLTXD_delay;
wire [0:31] DMA2LLTXD_delay;
wire [0:31] DMA3LLTXD_delay;
wire [0:31] PPCDMDCRDBUSOUT_delay;
wire [0:31] PPCDSDCRDBUSIN_delay;
wire [0:31] PPCMPLBABUS_delay;
wire [0:35] MIMCADDRESS_delay;
wire [0:3] APUFCMDECUDI_delay;
wire [0:3] APUFCMLOADBYTEADDR_delay;
wire [0:3] DMA0LLTXREM_delay;
wire [0:3] DMA1LLTXREM_delay;
wire [0:3] DMA2LLTXREM_delay;
wire [0:3] DMA3LLTXREM_delay;
wire [0:3] PPCMPLBSIZE_delay;
wire [0:3] PPCS0PLBMBUSY_delay;
wire [0:3] PPCS0PLBMIRQ_delay;
wire [0:3] PPCS0PLBMRDERR_delay;
wire [0:3] PPCS0PLBMWRERR_delay;
wire [0:3] PPCS0PLBRDWDADDR_delay;
wire [0:3] PPCS1PLBMBUSY_delay;
wire [0:3] PPCS1PLBMIRQ_delay;
wire [0:3] PPCS1PLBMRDERR_delay;
wire [0:3] PPCS1PLBMWRERR_delay;
wire [0:3] PPCS1PLBRDWDADDR_delay;
wire [0:4] C440TRCEXECUTIONSTATUS_delay;
wire [0:6] C440TRCTRACESTATUS_delay;
wire [0:7] C440DBGSYSTEMCONTROL_delay;
wire [0:9] PPCDMDCRABUS_delay;
wire [20:21] PPCDMDCRUABUS_delay;
wire [28:31] PPCMPLBUABUS_delay;

wire CPMC440CLKEN_delay;
wire CPMC440CLK_delay;
wire CPMC440CORECLOCKINACTIVE_delay;
wire CPMC440TIMERCLOCK_delay;
wire CPMDCRCLK_delay;
wire CPMDMA0LLCLK_delay;
wire CPMDMA1LLCLK_delay;
wire CPMDMA2LLCLK_delay;
wire CPMDMA3LLCLK_delay;
wire CPMFCMCLK_delay;
wire CPMINTERCONNECTCLKEN_delay;
wire CPMINTERCONNECTCLKNTO1_delay;
wire CPMINTERCONNECTCLK_delay;
wire CPMMCCLK_delay;
wire CPMPPCMPLBCLK_delay;
wire CPMPPCS0PLBCLK_delay;
wire CPMPPCS1PLBCLK_delay;
wire DBGC440DEBUGHALT_delay;
wire DBGC440UNCONDDEBUGEVENT_delay;
wire DCRPPCDMACK_delay;
wire DCRPPCDMTIMEOUTWAIT_delay;
wire DCRPPCDSREAD_delay;
wire DCRPPCDSWRITE_delay;
wire EICC440CRITIRQ_delay;
wire EICC440EXTIRQ_delay;
wire FCMAPUCONFIRMINSTR_delay;
wire FCMAPUDONE_delay;
wire FCMAPUEXCEPTION_delay;
wire FCMAPUFPSCRFEX_delay;
wire FCMAPURESULTVALID_delay;
wire FCMAPUSLEEPNOTREADY_delay;
wire JTGC440TCK_delay;
wire JTGC440TDI_delay;
wire JTGC440TMS_delay;
wire JTGC440TRSTNEG_delay;
wire LLDMA0RSTENGINEREQ_delay;
wire LLDMA0RXEOFN_delay;
wire LLDMA0RXEOPN_delay;
wire LLDMA0RXSOFN_delay;
wire LLDMA0RXSOPN_delay;
wire LLDMA0RXSRCRDYN_delay;
wire LLDMA0TXDSTRDYN_delay;
wire LLDMA1RSTENGINEREQ_delay;
wire LLDMA1RXEOFN_delay;
wire LLDMA1RXEOPN_delay;
wire LLDMA1RXSOFN_delay;
wire LLDMA1RXSOPN_delay;
wire LLDMA1RXSRCRDYN_delay;
wire LLDMA1TXDSTRDYN_delay;
wire LLDMA2RSTENGINEREQ_delay;
wire LLDMA2RXEOFN_delay;
wire LLDMA2RXEOPN_delay;
wire LLDMA2RXSOFN_delay;
wire LLDMA2RXSOPN_delay;
wire LLDMA2RXSRCRDYN_delay;
wire LLDMA2TXDSTRDYN_delay;
wire LLDMA3RSTENGINEREQ_delay;
wire LLDMA3RXEOFN_delay;
wire LLDMA3RXEOPN_delay;
wire LLDMA3RXSOFN_delay;
wire LLDMA3RXSOPN_delay;
wire LLDMA3RXSRCRDYN_delay;
wire LLDMA3TXDSTRDYN_delay;
wire MCMIADDRREADYTOACCEPT_delay;
wire MCMIREADDATAERR_delay;
wire MCMIREADDATAVALID_delay;
wire PLBPPCMADDRACK_delay;
wire PLBPPCMMBUSY_delay;
wire PLBPPCMMIRQ_delay;
wire PLBPPCMMRDERR_delay;
wire PLBPPCMMWRERR_delay;
wire PLBPPCMRDBTERM_delay;
wire PLBPPCMRDDACK_delay;
wire PLBPPCMRDPENDREQ_delay;
wire PLBPPCMREARBITRATE_delay;
wire PLBPPCMTIMEOUT_delay;
wire PLBPPCMWRBTERM_delay;
wire PLBPPCMWRDACK_delay;
wire PLBPPCMWRPENDREQ_delay;
wire PLBPPCS0ABORT_delay;
wire PLBPPCS0BUSLOCK_delay;
wire PLBPPCS0LOCKERR_delay;
wire PLBPPCS0PAVALID_delay;
wire PLBPPCS0RDBURST_delay;
wire PLBPPCS0RDPENDREQ_delay;
wire PLBPPCS0RDPRIM_delay;
wire PLBPPCS0RNW_delay;
wire PLBPPCS0SAVALID_delay;
wire PLBPPCS0WRBURST_delay;
wire PLBPPCS0WRPENDREQ_delay;
wire PLBPPCS0WRPRIM_delay;
wire PLBPPCS1ABORT_delay;
wire PLBPPCS1BUSLOCK_delay;
wire PLBPPCS1LOCKERR_delay;
wire PLBPPCS1PAVALID_delay;
wire PLBPPCS1RDBURST_delay;
wire PLBPPCS1RDPENDREQ_delay;
wire PLBPPCS1RDPRIM_delay;
wire PLBPPCS1RNW_delay;
wire PLBPPCS1SAVALID_delay;
wire PLBPPCS1WRBURST_delay;
wire PLBPPCS1WRPENDREQ_delay;
wire PLBPPCS1WRPRIM_delay;
wire RSTC440RESETCHIP_delay;
wire RSTC440RESETCORE_delay;
wire RSTC440RESETSYSTEM_delay;
wire TIEC440ENDIANRESET_delay;
wire TRCC440TRACEDISABLE_delay;
wire TRCC440TRIGGEREVENTIN_delay;
wire [0:127] FCMAPUSTOREDATA_delay;
wire [0:127] MCMIREADDATA_delay;
wire [0:127] PLBPPCMRDDBUS_delay;
wire [0:127] PLBPPCS0WRDBUS_delay;
wire [0:127] PLBPPCS1WRDBUS_delay;
wire [0:15] PLBPPCS0BE_delay;
wire [0:15] PLBPPCS0TATTRIBUTE_delay;
wire [0:15] PLBPPCS1BE_delay;
wire [0:15] PLBPPCS1TATTRIBUTE_delay;
wire [0:1] PLBPPCMRDPENDPRI_delay;
wire [0:1] PLBPPCMREQPRI_delay;
wire [0:1] PLBPPCMSSIZE_delay;
wire [0:1] PLBPPCMWRPENDPRI_delay;
wire [0:1] PLBPPCS0MASTERID_delay;
wire [0:1] PLBPPCS0MSIZE_delay;
wire [0:1] PLBPPCS0RDPENDPRI_delay;
wire [0:1] PLBPPCS0REQPRI_delay;
wire [0:1] PLBPPCS0WRPENDPRI_delay;
wire [0:1] PLBPPCS1MASTERID_delay;
wire [0:1] PLBPPCS1MSIZE_delay;
wire [0:1] PLBPPCS1RDPENDPRI_delay;
wire [0:1] PLBPPCS1REQPRI_delay;
wire [0:1] PLBPPCS1WRPENDPRI_delay;
wire [0:1] TIEC440DCURDLDCACHEPLBPRIO_delay;
wire [0:1] TIEC440DCURDNONCACHEPLBPRIO_delay;
wire [0:1] TIEC440DCURDTOUCHPLBPRIO_delay;
wire [0:1] TIEC440DCURDURGENTPLBPRIO_delay;
wire [0:1] TIEC440DCUWRFLUSHPLBPRIO_delay;
wire [0:1] TIEC440DCUWRSTOREPLBPRIO_delay;
wire [0:1] TIEC440DCUWRURGENTPLBPRIO_delay;
wire [0:1] TIEC440ICURDFETCHPLBPRIO_delay;
wire [0:1] TIEC440ICURDSPECPLBPRIO_delay;
wire [0:1] TIEC440ICURDTOUCHPLBPRIO_delay;
wire [0:1] TIEDCRBASEADDR_delay;
wire [0:2] PLBPPCS0TYPE_delay;
wire [0:2] PLBPPCS1TYPE_delay;
wire [0:31] DCRPPCDMDBUSIN_delay;
wire [0:31] DCRPPCDSDBUSOUT_delay;
wire [0:31] FCMAPURESULT_delay;
wire [0:31] LLDMA0RXD_delay;
wire [0:31] LLDMA1RXD_delay;
wire [0:31] LLDMA2RXD_delay;
wire [0:31] LLDMA3RXD_delay;
wire [0:31] PLBPPCS0ABUS_delay;
wire [0:31] PLBPPCS1ABUS_delay;
wire [0:3] FCMAPUCR_delay;
wire [0:3] LLDMA0RXREM_delay;
wire [0:3] LLDMA1RXREM_delay;
wire [0:3] LLDMA2RXREM_delay;
wire [0:3] LLDMA3RXREM_delay;
wire [0:3] PLBPPCMRDWDADDR_delay;
wire [0:3] PLBPPCS0SIZE_delay;
wire [0:3] PLBPPCS1SIZE_delay;
wire [0:3] TIEC440ERPNRESET_delay;
wire [0:3] TIEC440USERRESET_delay;
wire [0:4] DBGC440SYSTEMSTATUS_delay;
wire [0:9] DCRPPCDSABUS_delay;
wire [28:31] PLBPPCS0UABUS_delay;
wire [28:31] PLBPPCS1UABUS_delay;
wire [28:31] TIEC440PIR_delay;
wire [28:31] TIEC440PVR_delay;


assign #(out_delay) APUFCMDECFPUOP_OUT = APUFCMDECFPUOP_delay;
assign #(out_delay) APUFCMDECLDSTXFERSIZE_OUT = APUFCMDECLDSTXFERSIZE_delay;
assign #(out_delay) APUFCMDECLOAD_OUT = APUFCMDECLOAD_delay;
assign #(out_delay) APUFCMDECNONAUTON_OUT = APUFCMDECNONAUTON_delay;
assign #(out_delay) APUFCMDECSTORE_OUT = APUFCMDECSTORE_delay;
assign #(out_delay) APUFCMDECUDIVALID_OUT = APUFCMDECUDIVALID_delay;
assign #(out_delay) APUFCMDECUDI_OUT = APUFCMDECUDI_delay;
assign #(out_delay) APUFCMENDIAN_OUT = APUFCMENDIAN_delay;
assign #(out_delay) APUFCMFLUSH_OUT = APUFCMFLUSH_delay;
assign #(out_delay) APUFCMINSTRUCTION_OUT = APUFCMINSTRUCTION_delay;
assign #(out_delay) APUFCMINSTRVALID_OUT = APUFCMINSTRVALID_delay;
assign #(out_delay) APUFCMLOADBYTEADDR_OUT = APUFCMLOADBYTEADDR_delay;
assign #(out_delay) APUFCMLOADDATA_OUT = APUFCMLOADDATA_delay;
assign #(out_delay) APUFCMLOADDVALID_OUT = APUFCMLOADDVALID_delay;
assign #(out_delay) APUFCMMSRFE0_OUT = APUFCMMSRFE0_delay;
assign #(out_delay) APUFCMMSRFE1_OUT = APUFCMMSRFE1_delay;
assign #(out_delay) APUFCMNEXTINSTRREADY_OUT = APUFCMNEXTINSTRREADY_delay;
assign #(out_delay) APUFCMOPERANDVALID_OUT = APUFCMOPERANDVALID_delay;
assign #(out_delay) APUFCMRADATA_OUT = APUFCMRADATA_delay;
assign #(out_delay) APUFCMRBDATA_OUT = APUFCMRBDATA_delay;
assign #(out_delay) APUFCMWRITEBACKOK_OUT = APUFCMWRITEBACKOK_delay;
assign #(out_delay) C440CPMCORESLEEPREQ_OUT = C440CPMCORESLEEPREQ_delay;
assign #(out_delay) C440CPMDECIRPTREQ_OUT = C440CPMDECIRPTREQ_delay;
assign #(out_delay) C440CPMFITIRPTREQ_OUT = C440CPMFITIRPTREQ_delay;
assign #(out_delay) C440CPMMSRCE_OUT = C440CPMMSRCE_delay;
assign #(out_delay) C440CPMMSREE_OUT = C440CPMMSREE_delay;
assign #(out_delay) C440CPMTIMERRESETREQ_OUT = C440CPMTIMERRESETREQ_delay;
assign #(out_delay) C440CPMWDIRPTREQ_OUT = C440CPMWDIRPTREQ_delay;
assign #(out_delay) C440DBGSYSTEMCONTROL_OUT = C440DBGSYSTEMCONTROL_delay;
assign #(out_delay) C440JTGTDOEN_OUT = C440JTGTDOEN_delay;
assign #(out_delay) C440JTGTDO_OUT = C440JTGTDO_delay;
assign #(out_delay) C440MACHINECHECK_OUT = C440MACHINECHECK_delay;
assign #(out_delay) C440RSTCHIPRESETREQ_OUT = C440RSTCHIPRESETREQ_delay;
assign #(out_delay) C440RSTCORERESETREQ_OUT = C440RSTCORERESETREQ_delay;
assign #(out_delay) C440RSTSYSTEMRESETREQ_OUT = C440RSTSYSTEMRESETREQ_delay;
assign #(out_delay) C440TRCBRANCHSTATUS_OUT = C440TRCBRANCHSTATUS_delay;
assign #(out_delay) C440TRCCYCLE_OUT = C440TRCCYCLE_delay;
assign #(out_delay) C440TRCEXECUTIONSTATUS_OUT = C440TRCEXECUTIONSTATUS_delay;
assign #(out_delay) C440TRCTRACESTATUS_OUT = C440TRCTRACESTATUS_delay;
assign #(out_delay) C440TRCTRIGGEREVENTOUT_OUT = C440TRCTRIGGEREVENTOUT_delay;
assign #(out_delay) C440TRCTRIGGEREVENTTYPE_OUT = C440TRCTRIGGEREVENTTYPE_delay;
assign #(out_delay) DMA0LLRSTENGINEACK_OUT = DMA0LLRSTENGINEACK_delay;
assign #(out_delay) DMA0LLRXDSTRDYN_OUT = DMA0LLRXDSTRDYN_delay;
assign #(out_delay) DMA0LLTXD_OUT = DMA0LLTXD_delay;
assign #(out_delay) DMA0LLTXEOFN_OUT = DMA0LLTXEOFN_delay;
assign #(out_delay) DMA0LLTXEOPN_OUT = DMA0LLTXEOPN_delay;
assign #(out_delay) DMA0LLTXREM_OUT = DMA0LLTXREM_delay;
assign #(out_delay) DMA0LLTXSOFN_OUT = DMA0LLTXSOFN_delay;
assign #(out_delay) DMA0LLTXSOPN_OUT = DMA0LLTXSOPN_delay;
assign #(out_delay) DMA0LLTXSRCRDYN_OUT = DMA0LLTXSRCRDYN_delay;
assign #(out_delay) DMA0RXIRQ_OUT = DMA0RXIRQ_delay;
assign #(out_delay) DMA0TXIRQ_OUT = DMA0TXIRQ_delay;
assign #(out_delay) DMA1LLRSTENGINEACK_OUT = DMA1LLRSTENGINEACK_delay;
assign #(out_delay) DMA1LLRXDSTRDYN_OUT = DMA1LLRXDSTRDYN_delay;
assign #(out_delay) DMA1LLTXD_OUT = DMA1LLTXD_delay;
assign #(out_delay) DMA1LLTXEOFN_OUT = DMA1LLTXEOFN_delay;
assign #(out_delay) DMA1LLTXEOPN_OUT = DMA1LLTXEOPN_delay;
assign #(out_delay) DMA1LLTXREM_OUT = DMA1LLTXREM_delay;
assign #(out_delay) DMA1LLTXSOFN_OUT = DMA1LLTXSOFN_delay;
assign #(out_delay) DMA1LLTXSOPN_OUT = DMA1LLTXSOPN_delay;
assign #(out_delay) DMA1LLTXSRCRDYN_OUT = DMA1LLTXSRCRDYN_delay;
assign #(out_delay) DMA1RXIRQ_OUT = DMA1RXIRQ_delay;
assign #(out_delay) DMA1TXIRQ_OUT = DMA1TXIRQ_delay;
assign #(out_delay) DMA2LLRSTENGINEACK_OUT = DMA2LLRSTENGINEACK_delay;
assign #(out_delay) DMA2LLRXDSTRDYN_OUT = DMA2LLRXDSTRDYN_delay;
assign #(out_delay) DMA2LLTXD_OUT = DMA2LLTXD_delay;
assign #(out_delay) DMA2LLTXEOFN_OUT = DMA2LLTXEOFN_delay;
assign #(out_delay) DMA2LLTXEOPN_OUT = DMA2LLTXEOPN_delay;
assign #(out_delay) DMA2LLTXREM_OUT = DMA2LLTXREM_delay;
assign #(out_delay) DMA2LLTXSOFN_OUT = DMA2LLTXSOFN_delay;
assign #(out_delay) DMA2LLTXSOPN_OUT = DMA2LLTXSOPN_delay;
assign #(out_delay) DMA2LLTXSRCRDYN_OUT = DMA2LLTXSRCRDYN_delay;
assign #(out_delay) DMA2RXIRQ_OUT = DMA2RXIRQ_delay;
assign #(out_delay) DMA2TXIRQ_OUT = DMA2TXIRQ_delay;
assign #(out_delay) DMA3LLRSTENGINEACK_OUT = DMA3LLRSTENGINEACK_delay;
assign #(out_delay) DMA3LLRXDSTRDYN_OUT = DMA3LLRXDSTRDYN_delay;
assign #(out_delay) DMA3LLTXD_OUT = DMA3LLTXD_delay;
assign #(out_delay) DMA3LLTXEOFN_OUT = DMA3LLTXEOFN_delay;
assign #(out_delay) DMA3LLTXEOPN_OUT = DMA3LLTXEOPN_delay;
assign #(out_delay) DMA3LLTXREM_OUT = DMA3LLTXREM_delay;
assign #(out_delay) DMA3LLTXSOFN_OUT = DMA3LLTXSOFN_delay;
assign #(out_delay) DMA3LLTXSOPN_OUT = DMA3LLTXSOPN_delay;
assign #(out_delay) DMA3LLTXSRCRDYN_OUT = DMA3LLTXSRCRDYN_delay;
assign #(out_delay) DMA3RXIRQ_OUT = DMA3RXIRQ_delay;
assign #(out_delay) DMA3TXIRQ_OUT = DMA3TXIRQ_delay;
assign #(out_delay) MIMCADDRESSVALID_OUT = MIMCADDRESSVALID_delay;
assign #(out_delay) MIMCADDRESS_OUT = MIMCADDRESS_delay;
assign #(out_delay) MIMCBANKCONFLICT_OUT = MIMCBANKCONFLICT_delay;
assign #(out_delay) MIMCBYTEENABLE_OUT = MIMCBYTEENABLE_delay;
assign #(out_delay) MIMCREADNOTWRITE_OUT = MIMCREADNOTWRITE_delay;
assign #(out_delay) MIMCROWCONFLICT_OUT = MIMCROWCONFLICT_delay;
assign #(out_delay) MIMCWRITEDATAVALID_OUT = MIMCWRITEDATAVALID_delay;
assign #(out_delay) MIMCWRITEDATA_OUT = MIMCWRITEDATA_delay;
assign #(out_delay) PPCCPMINTERCONNECTBUSY_OUT = PPCCPMINTERCONNECTBUSY_delay;
assign #(out_delay) PPCDMDCRABUS_OUT = PPCDMDCRABUS_delay;
assign #(out_delay) PPCDMDCRDBUSOUT_OUT = PPCDMDCRDBUSOUT_delay;
assign #(out_delay) PPCDMDCRREAD_OUT = PPCDMDCRREAD_delay;
assign #(out_delay) PPCDMDCRUABUS_OUT = PPCDMDCRUABUS_delay;
assign #(out_delay) PPCDMDCRWRITE_OUT = PPCDMDCRWRITE_delay;
assign #(out_delay) PPCDSDCRACK_OUT = PPCDSDCRACK_delay;
assign #(out_delay) PPCDSDCRDBUSIN_OUT = PPCDSDCRDBUSIN_delay;
assign #(out_delay) PPCDSDCRTIMEOUTWAIT_OUT = PPCDSDCRTIMEOUTWAIT_delay;
assign #(out_delay) PPCEICINTERCONNECTIRQ_OUT = PPCEICINTERCONNECTIRQ_delay;
assign #(out_delay) PPCMPLBABORT_OUT = PPCMPLBABORT_delay;
assign #(out_delay) PPCMPLBABUS_OUT = PPCMPLBABUS_delay;
assign #(out_delay) PPCMPLBBE_OUT = PPCMPLBBE_delay;
assign #(out_delay) PPCMPLBBUSLOCK_OUT = PPCMPLBBUSLOCK_delay;
assign #(out_delay) PPCMPLBLOCKERR_OUT = PPCMPLBLOCKERR_delay;
assign #(out_delay) PPCMPLBPRIORITY_OUT = PPCMPLBPRIORITY_delay;
assign #(out_delay) PPCMPLBRDBURST_OUT = PPCMPLBRDBURST_delay;
assign #(out_delay) PPCMPLBREQUEST_OUT = PPCMPLBREQUEST_delay;
assign #(out_delay) PPCMPLBRNW_OUT = PPCMPLBRNW_delay;
assign #(out_delay) PPCMPLBSIZE_OUT = PPCMPLBSIZE_delay;
assign #(out_delay) PPCMPLBTATTRIBUTE_OUT = PPCMPLBTATTRIBUTE_delay;
assign #(out_delay) PPCMPLBTYPE_OUT = PPCMPLBTYPE_delay;
assign #(out_delay) PPCMPLBUABUS_OUT = PPCMPLBUABUS_delay;
assign #(out_delay) PPCMPLBWRBURST_OUT = PPCMPLBWRBURST_delay;
assign #(out_delay) PPCMPLBWRDBUS_OUT = PPCMPLBWRDBUS_delay;
assign #(out_delay) PPCS0PLBADDRACK_OUT = PPCS0PLBADDRACK_delay;
assign #(out_delay) PPCS0PLBMBUSY_OUT = PPCS0PLBMBUSY_delay;
assign #(out_delay) PPCS0PLBMIRQ_OUT = PPCS0PLBMIRQ_delay;
assign #(out_delay) PPCS0PLBMRDERR_OUT = PPCS0PLBMRDERR_delay;
assign #(out_delay) PPCS0PLBMWRERR_OUT = PPCS0PLBMWRERR_delay;
assign #(out_delay) PPCS0PLBRDBTERM_OUT = PPCS0PLBRDBTERM_delay;
assign #(out_delay) PPCS0PLBRDCOMP_OUT = PPCS0PLBRDCOMP_delay;
assign #(out_delay) PPCS0PLBRDDACK_OUT = PPCS0PLBRDDACK_delay;
assign #(out_delay) PPCS0PLBRDDBUS_OUT = PPCS0PLBRDDBUS_delay;
assign #(out_delay) PPCS0PLBRDWDADDR_OUT = PPCS0PLBRDWDADDR_delay;
assign #(out_delay) PPCS0PLBREARBITRATE_OUT = PPCS0PLBREARBITRATE_delay;
assign #(out_delay) PPCS0PLBSSIZE_OUT = PPCS0PLBSSIZE_delay;
assign #(out_delay) PPCS0PLBWAIT_OUT = PPCS0PLBWAIT_delay;
assign #(out_delay) PPCS0PLBWRBTERM_OUT = PPCS0PLBWRBTERM_delay;
assign #(out_delay) PPCS0PLBWRCOMP_OUT = PPCS0PLBWRCOMP_delay;
assign #(out_delay) PPCS0PLBWRDACK_OUT = PPCS0PLBWRDACK_delay;
assign #(out_delay) PPCS1PLBADDRACK_OUT = PPCS1PLBADDRACK_delay;
assign #(out_delay) PPCS1PLBMBUSY_OUT = PPCS1PLBMBUSY_delay;
assign #(out_delay) PPCS1PLBMIRQ_OUT = PPCS1PLBMIRQ_delay;
assign #(out_delay) PPCS1PLBMRDERR_OUT = PPCS1PLBMRDERR_delay;
assign #(out_delay) PPCS1PLBMWRERR_OUT = PPCS1PLBMWRERR_delay;
assign #(out_delay) PPCS1PLBRDBTERM_OUT = PPCS1PLBRDBTERM_delay;
assign #(out_delay) PPCS1PLBRDCOMP_OUT = PPCS1PLBRDCOMP_delay;
assign #(out_delay) PPCS1PLBRDDACK_OUT = PPCS1PLBRDDACK_delay;
assign #(out_delay) PPCS1PLBRDDBUS_OUT = PPCS1PLBRDDBUS_delay;
assign #(out_delay) PPCS1PLBRDWDADDR_OUT = PPCS1PLBRDWDADDR_delay;
assign #(out_delay) PPCS1PLBREARBITRATE_OUT = PPCS1PLBREARBITRATE_delay;
assign #(out_delay) PPCS1PLBSSIZE_OUT = PPCS1PLBSSIZE_delay;
assign #(out_delay) PPCS1PLBWAIT_OUT = PPCS1PLBWAIT_delay;
assign #(out_delay) PPCS1PLBWRBTERM_OUT = PPCS1PLBWRBTERM_delay;
assign #(out_delay) PPCS1PLBWRCOMP_OUT = PPCS1PLBWRCOMP_delay;
assign #(out_delay) PPCS1PLBWRDACK_OUT = PPCS1PLBWRDACK_delay;

// assign #(CLK_DELAY) CPMC440CLK_delay = CPMC440CLK_IN;
assign #(CLK_DELAY) CPMC440TIMERCLOCK_delay = CPMC440TIMERCLOCK_IN;
// assign #(CLK_DELAY) CPMDCRCLK_delay = CPMDCRCLK_IN;
// assign #(CLK_DELAY) CPMDMA0LLCLK_delay = CPMDMA0LLCLK_IN;
// assign #(CLK_DELAY) CPMDMA1LLCLK_delay = CPMDMA1LLCLK_IN;
// assign #(CLK_DELAY) CPMDMA2LLCLK_delay = CPMDMA2LLCLK_IN;
// assign #(CLK_DELAY) CPMDMA3LLCLK_delay = CPMDMA3LLCLK_IN;
// assign #(CLK_DELAY) CPMFCMCLK_delay = CPMFCMCLK_IN;
// assign #(CLK_DELAY) CPMINTERCONNECTCLK_delay = CPMINTERCONNECTCLK_IN;
// assign #(CLK_DELAY) CPMMCCLK_delay = CPMMCCLK_IN;
// assign #(CLK_DELAY) CPMPPCMPLBCLK_delay = CPMPPCMPLBCLK_IN;
// assign #(CLK_DELAY) CPMPPCS0PLBCLK_delay = CPMPPCS0PLBCLK_IN;
// assign #(CLK_DELAY) CPMPPCS1PLBCLK_delay = CPMPPCS1PLBCLK_IN;
// assign #(CLK_DELAY) JTGC440TCK_delay = JTGC440TCK_IN;

assign #(in_delay) CPMC440CLKEN_delay = CPMC440CLKEN_IN;
// assign #(in_delay) CPMC440CORECLOCKINACTIVE_delay = CPMC440CORECLOCKINACTIVE_IN;
assign #(in_delay) CPMINTERCONNECTCLKEN_delay = CPMINTERCONNECTCLKEN_IN;
// assign #(in_delay) CPMINTERCONNECTCLKNTO1_delay = CPMINTERCONNECTCLKNTO1_IN;
// assign #(in_delay) DBGC440DEBUGHALT_delay = DBGC440DEBUGHALT_IN;
// assign #(in_delay) DBGC440SYSTEMSTATUS_delay = DBGC440SYSTEMSTATUS_IN;
// assign #(in_delay) DBGC440UNCONDDEBUGEVENT_delay = DBGC440UNCONDDEBUGEVENT_IN;
// assign #(in_delay) DCRPPCDMACK_delay = DCRPPCDMACK_IN;
// assign #(in_delay) DCRPPCDMDBUSIN_delay = DCRPPCDMDBUSIN_IN;
// assign #(in_delay) DCRPPCDMTIMEOUTWAIT_delay = DCRPPCDMTIMEOUTWAIT_IN;
// assign #(in_delay) DCRPPCDSABUS_delay = DCRPPCDSABUS_IN;
// assign #(in_delay) DCRPPCDSDBUSOUT_delay = DCRPPCDSDBUSOUT_IN;
// assign #(in_delay) DCRPPCDSREAD_delay = DCRPPCDSREAD_IN;
// assign #(in_delay) DCRPPCDSWRITE_delay = DCRPPCDSWRITE_IN;
assign #(in_delay) EICC440CRITIRQ_delay = EICC440CRITIRQ_IN;
assign #(in_delay) EICC440EXTIRQ_delay = EICC440EXTIRQ_IN;
// assign #(in_delay) FCMAPUCONFIRMINSTR_delay = FCMAPUCONFIRMINSTR_IN;
// assign #(in_delay) FCMAPUCR_delay = FCMAPUCR_IN;
// assign #(in_delay) FCMAPUDONE_delay = FCMAPUDONE_IN;
// assign #(in_delay) FCMAPUEXCEPTION_delay = FCMAPUEXCEPTION_IN;
// assign #(in_delay) FCMAPUFPSCRFEX_delay = FCMAPUFPSCRFEX_IN;
// assign #(in_delay) FCMAPURESULTVALID_delay = FCMAPURESULTVALID_IN;
// assign #(in_delay) FCMAPURESULT_delay = FCMAPURESULT_IN;
// assign #(in_delay) FCMAPUSLEEPNOTREADY_delay = FCMAPUSLEEPNOTREADY_IN;
// assign #(in_delay) FCMAPUSTOREDATA_delay = FCMAPUSTOREDATA_IN;
// assign #(in_delay) JTGC440TDI_delay = JTGC440TDI_IN;
// assign #(in_delay) JTGC440TMS_delay = JTGC440TMS_IN;
assign #(in_delay) JTGC440TRSTNEG_delay = JTGC440TRSTNEG_IN;
// assign #(in_delay) LLDMA0RSTENGINEREQ_delay = LLDMA0RSTENGINEREQ_IN;
// assign #(in_delay) LLDMA0RXD_delay = LLDMA0RXD_IN;
// assign #(in_delay) LLDMA0RXEOFN_delay = LLDMA0RXEOFN_IN;
// assign #(in_delay) LLDMA0RXEOPN_delay = LLDMA0RXEOPN_IN;
// assign #(in_delay) LLDMA0RXREM_delay = LLDMA0RXREM_IN;
// assign #(in_delay) LLDMA0RXSOFN_delay = LLDMA0RXSOFN_IN;
// assign #(in_delay) LLDMA0RXSOPN_delay = LLDMA0RXSOPN_IN;
// assign #(in_delay) LLDMA0RXSRCRDYN_delay = LLDMA0RXSRCRDYN_IN;
// assign #(in_delay) LLDMA0TXDSTRDYN_delay = LLDMA0TXDSTRDYN_IN;
// assign #(in_delay) LLDMA1RSTENGINEREQ_delay = LLDMA1RSTENGINEREQ_IN;
// assign #(in_delay) LLDMA1RXD_delay = LLDMA1RXD_IN;
// assign #(in_delay) LLDMA1RXEOFN_delay = LLDMA1RXEOFN_IN;
// assign #(in_delay) LLDMA1RXEOPN_delay = LLDMA1RXEOPN_IN;
// assign #(in_delay) LLDMA1RXREM_delay = LLDMA1RXREM_IN;
// assign #(in_delay) LLDMA1RXSOFN_delay = LLDMA1RXSOFN_IN;
// assign #(in_delay) LLDMA1RXSOPN_delay = LLDMA1RXSOPN_IN;
// assign #(in_delay) LLDMA1RXSRCRDYN_delay = LLDMA1RXSRCRDYN_IN;
// assign #(in_delay) LLDMA1TXDSTRDYN_delay = LLDMA1TXDSTRDYN_IN;
// assign #(in_delay) LLDMA2RSTENGINEREQ_delay = LLDMA2RSTENGINEREQ_IN;
// assign #(in_delay) LLDMA2RXD_delay = LLDMA2RXD_IN;
// assign #(in_delay) LLDMA2RXEOFN_delay = LLDMA2RXEOFN_IN;
// assign #(in_delay) LLDMA2RXEOPN_delay = LLDMA2RXEOPN_IN;
// assign #(in_delay) LLDMA2RXREM_delay = LLDMA2RXREM_IN;
// assign #(in_delay) LLDMA2RXSOFN_delay = LLDMA2RXSOFN_IN;
// assign #(in_delay) LLDMA2RXSOPN_delay = LLDMA2RXSOPN_IN;
// assign #(in_delay) LLDMA2RXSRCRDYN_delay = LLDMA2RXSRCRDYN_IN;
// assign #(in_delay) LLDMA2TXDSTRDYN_delay = LLDMA2TXDSTRDYN_IN;
// assign #(in_delay) LLDMA3RSTENGINEREQ_delay = LLDMA3RSTENGINEREQ_IN;
// assign #(in_delay) LLDMA3RXD_delay = LLDMA3RXD_IN;
// assign #(in_delay) LLDMA3RXEOFN_delay = LLDMA3RXEOFN_IN;
// assign #(in_delay) LLDMA3RXEOPN_delay = LLDMA3RXEOPN_IN;
// assign #(in_delay) LLDMA3RXREM_delay = LLDMA3RXREM_IN;
// assign #(in_delay) LLDMA3RXSOFN_delay = LLDMA3RXSOFN_IN;
// assign #(in_delay) LLDMA3RXSOPN_delay = LLDMA3RXSOPN_IN;
// assign #(in_delay) LLDMA3RXSRCRDYN_delay = LLDMA3RXSRCRDYN_IN;
// assign #(in_delay) LLDMA3TXDSTRDYN_delay = LLDMA3TXDSTRDYN_IN;
// assign #(in_delay) MCMIADDRREADYTOACCEPT_delay = MCMIADDRREADYTOACCEPT_IN;
// assign #(in_delay) MCMIREADDATAERR_delay = MCMIREADDATAERR_IN;
// assign #(in_delay) MCMIREADDATAVALID_delay = MCMIREADDATAVALID_IN;
// assign #(in_delay) MCMIREADDATA_delay = MCMIREADDATA_IN;
// assign #(in_delay) PLBPPCMADDRACK_delay = PLBPPCMADDRACK_IN;
// assign #(in_delay) PLBPPCMMBUSY_delay = PLBPPCMMBUSY_IN;
// assign #(in_delay) PLBPPCMMIRQ_delay = PLBPPCMMIRQ_IN;
// assign #(in_delay) PLBPPCMMRDERR_delay = PLBPPCMMRDERR_IN;
// assign #(in_delay) PLBPPCMMWRERR_delay = PLBPPCMMWRERR_IN;
// assign #(in_delay) PLBPPCMRDBTERM_delay = PLBPPCMRDBTERM_IN;
// assign #(in_delay) PLBPPCMRDDACK_delay = PLBPPCMRDDACK_IN;
// assign #(in_delay) PLBPPCMRDDBUS_delay = PLBPPCMRDDBUS_IN;
// assign #(in_delay) PLBPPCMRDPENDPRI_delay = PLBPPCMRDPENDPRI_IN;
// assign #(in_delay) PLBPPCMRDPENDREQ_delay = PLBPPCMRDPENDREQ_IN;
// assign #(in_delay) PLBPPCMRDWDADDR_delay = PLBPPCMRDWDADDR_IN;
// assign #(in_delay) PLBPPCMREARBITRATE_delay = PLBPPCMREARBITRATE_IN;
// assign #(in_delay) PLBPPCMREQPRI_delay = PLBPPCMREQPRI_IN;
// assign #(in_delay) PLBPPCMSSIZE_delay = PLBPPCMSSIZE_IN;
// assign #(in_delay) PLBPPCMTIMEOUT_delay = PLBPPCMTIMEOUT_IN;
// assign #(in_delay) PLBPPCMWRBTERM_delay = PLBPPCMWRBTERM_IN;
// assign #(in_delay) PLBPPCMWRDACK_delay = PLBPPCMWRDACK_IN;
// assign #(in_delay) PLBPPCMWRPENDPRI_delay = PLBPPCMWRPENDPRI_IN;
// assign #(in_delay) PLBPPCMWRPENDREQ_delay = PLBPPCMWRPENDREQ_IN;
// assign #(in_delay) PLBPPCS0ABORT_delay = PLBPPCS0ABORT_IN;
// assign #(in_delay) PLBPPCS0ABUS_delay = PLBPPCS0ABUS_IN;
// assign #(in_delay) PLBPPCS0BE_delay = PLBPPCS0BE_IN;
// assign #(in_delay) PLBPPCS0BUSLOCK_delay = PLBPPCS0BUSLOCK_IN;
// assign #(in_delay) PLBPPCS0LOCKERR_delay = PLBPPCS0LOCKERR_IN;
// assign #(in_delay) PLBPPCS0MASTERID_delay = PLBPPCS0MASTERID_IN;
// assign #(in_delay) PLBPPCS0MSIZE_delay = PLBPPCS0MSIZE_IN;
// assign #(in_delay) PLBPPCS0PAVALID_delay = PLBPPCS0PAVALID_IN;
// assign #(in_delay) PLBPPCS0RDBURST_delay = PLBPPCS0RDBURST_IN;
// assign #(in_delay) PLBPPCS0RDPENDPRI_delay = PLBPPCS0RDPENDPRI_IN;
// assign #(in_delay) PLBPPCS0RDPENDREQ_delay = PLBPPCS0RDPENDREQ_IN;
// assign #(in_delay) PLBPPCS0RDPRIM_delay = PLBPPCS0RDPRIM_IN;
// assign #(in_delay) PLBPPCS0REQPRI_delay = PLBPPCS0REQPRI_IN;
// assign #(in_delay) PLBPPCS0RNW_delay = PLBPPCS0RNW_IN;
// assign #(in_delay) PLBPPCS0SAVALID_delay = PLBPPCS0SAVALID_IN;
// assign #(in_delay) PLBPPCS0SIZE_delay = PLBPPCS0SIZE_IN;
// assign #(in_delay) PLBPPCS0TATTRIBUTE_delay = PLBPPCS0TATTRIBUTE_IN;
// assign #(in_delay) PLBPPCS0TYPE_delay = PLBPPCS0TYPE_IN;
// assign #(in_delay) PLBPPCS0UABUS_delay = PLBPPCS0UABUS_IN;
// assign #(in_delay) PLBPPCS0WRBURST_delay = PLBPPCS0WRBURST_IN;
// assign #(in_delay) PLBPPCS0WRDBUS_delay = PLBPPCS0WRDBUS_IN;
// assign #(in_delay) PLBPPCS0WRPENDPRI_delay = PLBPPCS0WRPENDPRI_IN;
// assign #(in_delay) PLBPPCS0WRPENDREQ_delay = PLBPPCS0WRPENDREQ_IN;
// assign #(in_delay) PLBPPCS0WRPRIM_delay = PLBPPCS0WRPRIM_IN;
// assign #(in_delay) PLBPPCS1ABORT_delay = PLBPPCS1ABORT_IN;
// assign #(in_delay) PLBPPCS1ABUS_delay = PLBPPCS1ABUS_IN;
// assign #(in_delay) PLBPPCS1BE_delay = PLBPPCS1BE_IN;
// assign #(in_delay) PLBPPCS1BUSLOCK_delay = PLBPPCS1BUSLOCK_IN;
// assign #(in_delay) PLBPPCS1LOCKERR_delay = PLBPPCS1LOCKERR_IN;
// assign #(in_delay) PLBPPCS1MASTERID_delay = PLBPPCS1MASTERID_IN;
// assign #(in_delay) PLBPPCS1MSIZE_delay = PLBPPCS1MSIZE_IN;
// assign #(in_delay) PLBPPCS1PAVALID_delay = PLBPPCS1PAVALID_IN;
// assign #(in_delay) PLBPPCS1RDBURST_delay = PLBPPCS1RDBURST_IN;
// assign #(in_delay) PLBPPCS1RDPENDPRI_delay = PLBPPCS1RDPENDPRI_IN;
// assign #(in_delay) PLBPPCS1RDPENDREQ_delay = PLBPPCS1RDPENDREQ_IN;
// assign #(in_delay) PLBPPCS1RDPRIM_delay = PLBPPCS1RDPRIM_IN;
// assign #(in_delay) PLBPPCS1REQPRI_delay = PLBPPCS1REQPRI_IN;
// assign #(in_delay) PLBPPCS1RNW_delay = PLBPPCS1RNW_IN;
// assign #(in_delay) PLBPPCS1SAVALID_delay = PLBPPCS1SAVALID_IN;
// assign #(in_delay) PLBPPCS1SIZE_delay = PLBPPCS1SIZE_IN;
// assign #(in_delay) PLBPPCS1TATTRIBUTE_delay = PLBPPCS1TATTRIBUTE_IN;
// assign #(in_delay) PLBPPCS1TYPE_delay = PLBPPCS1TYPE_IN;
// assign #(in_delay) PLBPPCS1UABUS_delay = PLBPPCS1UABUS_IN;
// assign #(in_delay) PLBPPCS1WRBURST_delay = PLBPPCS1WRBURST_IN;
// assign #(in_delay) PLBPPCS1WRDBUS_delay = PLBPPCS1WRDBUS_IN;
// assign #(in_delay) PLBPPCS1WRPENDPRI_delay = PLBPPCS1WRPENDPRI_IN;
// assign #(in_delay) PLBPPCS1WRPENDREQ_delay = PLBPPCS1WRPENDREQ_IN;
// assign #(in_delay) PLBPPCS1WRPRIM_delay = PLBPPCS1WRPRIM_IN;
assign #(in_delay) RSTC440RESETCHIP_delay = RSTC440RESETCHIP_IN;
assign #(in_delay) RSTC440RESETCORE_delay = RSTC440RESETCORE_IN;
assign #(in_delay) RSTC440RESETSYSTEM_delay = RSTC440RESETSYSTEM_IN;
assign #(in_delay) TIEC440DCURDLDCACHEPLBPRIO_delay = TIEC440DCURDLDCACHEPLBPRIO_IN;
assign #(in_delay) TIEC440DCURDNONCACHEPLBPRIO_delay = TIEC440DCURDNONCACHEPLBPRIO_IN;
assign #(in_delay) TIEC440DCURDTOUCHPLBPRIO_delay = TIEC440DCURDTOUCHPLBPRIO_IN;
assign #(in_delay) TIEC440DCURDURGENTPLBPRIO_delay = TIEC440DCURDURGENTPLBPRIO_IN;
assign #(in_delay) TIEC440DCUWRFLUSHPLBPRIO_delay = TIEC440DCUWRFLUSHPLBPRIO_IN;
assign #(in_delay) TIEC440DCUWRSTOREPLBPRIO_delay = TIEC440DCUWRSTOREPLBPRIO_IN;
assign #(in_delay) TIEC440DCUWRURGENTPLBPRIO_delay = TIEC440DCUWRURGENTPLBPRIO_IN;
assign #(in_delay) TIEC440ENDIANRESET_delay = TIEC440ENDIANRESET_IN;
assign #(in_delay) TIEC440ERPNRESET_delay = TIEC440ERPNRESET_IN;
assign #(in_delay) TIEC440ICURDFETCHPLBPRIO_delay = TIEC440ICURDFETCHPLBPRIO_IN;
assign #(in_delay) TIEC440ICURDSPECPLBPRIO_delay = TIEC440ICURDSPECPLBPRIO_IN;
assign #(in_delay) TIEC440ICURDTOUCHPLBPRIO_delay = TIEC440ICURDTOUCHPLBPRIO_IN;
assign #(in_delay) TIEC440PIR_delay = TIEC440PIR_IN;
assign #(in_delay) TIEC440PVR_delay = TIEC440PVR_IN;
assign #(in_delay) TIEC440USERRESET_delay = TIEC440USERRESET_IN;
assign #(in_delay) TIEDCRBASEADDR_delay = TIEDCRBASEADDR_IN;
// assign #(in_delay) TRCC440TRACEDISABLE_delay = TRCC440TRACEDISABLE_IN;
// assign #(in_delay) TRCC440TRIGGEREVENTIN_delay = TRCC440TRIGGEREVENTIN_IN;


PPC440_SWIFT ppc440_swift_1 (
	.APU_CONTROL (APU_CONTROL),
	.APU_UDI0 (APU_UDI0),
	.APU_UDI1 (APU_UDI1),
	.APU_UDI10 (APU_UDI10),
	.APU_UDI11 (APU_UDI11),
	.APU_UDI12 (APU_UDI12),
	.APU_UDI13 (APU_UDI13),
	.APU_UDI14 (APU_UDI14),
	.APU_UDI15 (APU_UDI15),
	.APU_UDI2 (APU_UDI2),
	.APU_UDI3 (APU_UDI3),
	.APU_UDI4 (APU_UDI4),
	.APU_UDI5 (APU_UDI5),
	.APU_UDI6 (APU_UDI6),
	.APU_UDI7 (APU_UDI7),
	.APU_UDI8 (APU_UDI8),
	.APU_UDI9 (APU_UDI9),
	.CLOCK_DELAY (CLOCK_DELAY_BINARY),
	.DCR_AUTOLOCK_ENABLE (DCR_AUTOLOCK_ENABLE_BINARY),
	.DMA0_CONTROL (DMA0_CONTROL),
	.DMA0_RXCHANNELCTRL (DMA0_RXCHANNELCTRL),
	.DMA0_RXIRQTIMER (DMA0_RXIRQTIMER),
	.DMA0_TXCHANNELCTRL (DMA0_TXCHANNELCTRL),
	.DMA0_TXIRQTIMER (DMA0_TXIRQTIMER),
	.DMA1_CONTROL (DMA1_CONTROL),
	.DMA1_RXCHANNELCTRL (DMA1_RXCHANNELCTRL),
	.DMA1_RXIRQTIMER (DMA1_RXIRQTIMER),
	.DMA1_TXCHANNELCTRL (DMA1_TXCHANNELCTRL),
	.DMA1_TXIRQTIMER (DMA1_TXIRQTIMER),
	.DMA2_CONTROL (DMA2_CONTROL),
	.DMA2_RXCHANNELCTRL (DMA2_RXCHANNELCTRL),
	.DMA2_RXIRQTIMER (DMA2_RXIRQTIMER),
	.DMA2_TXCHANNELCTRL (DMA2_TXCHANNELCTRL),
	.DMA2_TXIRQTIMER (DMA2_TXIRQTIMER),
	.DMA3_CONTROL (DMA3_CONTROL),
	.DMA3_RXCHANNELCTRL (DMA3_RXCHANNELCTRL),
	.DMA3_RXIRQTIMER (DMA3_RXIRQTIMER),
	.DMA3_TXCHANNELCTRL (DMA3_TXCHANNELCTRL),
	.DMA3_TXIRQTIMER (DMA3_TXIRQTIMER),
	.INTERCONNECT_IMASK (INTERCONNECT_IMASK),
	.INTERCONNECT_TMPL_SEL (INTERCONNECT_TMPL_SEL),
	.MI_ARBCONFIG (MI_ARBCONFIG),
	.MI_BANKCONFLICT_MASK (MI_BANKCONFLICT_MASK),
	.MI_CONTROL (MI_CONTROL),
	.MI_ROWCONFLICT_MASK (MI_ROWCONFLICT_MASK),
	.PPCDM_ASYNCMODE (PPCDM_ASYNCMODE_BINARY),
	.PPCDS_ASYNCMODE (PPCDS_ASYNCMODE_BINARY),
	.PPCM_ARBCONFIG (PPCM_ARBCONFIG),
	.PPCM_CONTROL (PPCM_CONTROL),
	.PPCM_COUNTER (PPCM_COUNTER),
	.PPCS0_ADDRMAP_TMPL0 (PPCS0_ADDRMAP_TMPL0),
	.PPCS0_ADDRMAP_TMPL1 (PPCS0_ADDRMAP_TMPL1),
	.PPCS0_ADDRMAP_TMPL2 (PPCS0_ADDRMAP_TMPL2),
	.PPCS0_ADDRMAP_TMPL3 (PPCS0_ADDRMAP_TMPL3),
	.PPCS0_CONTROL (PPCS0_CONTROL),
	.PPCS0_WIDTH_128N64 (PPCS0_WIDTH_128N64_BINARY),
	.PPCS1_ADDRMAP_TMPL0 (PPCS1_ADDRMAP_TMPL0),
	.PPCS1_ADDRMAP_TMPL1 (PPCS1_ADDRMAP_TMPL1),
	.PPCS1_ADDRMAP_TMPL2 (PPCS1_ADDRMAP_TMPL2),
	.PPCS1_ADDRMAP_TMPL3 (PPCS1_ADDRMAP_TMPL3),
	.PPCS1_CONTROL (PPCS1_CONTROL),
	.PPCS1_WIDTH_128N64 (PPCS1_WIDTH_128N64_BINARY),
	.XBAR_ADDRMAP_TMPL0 (XBAR_ADDRMAP_TMPL0),
	.XBAR_ADDRMAP_TMPL1 (XBAR_ADDRMAP_TMPL1),
	.XBAR_ADDRMAP_TMPL2 (XBAR_ADDRMAP_TMPL2),
	.XBAR_ADDRMAP_TMPL3 (XBAR_ADDRMAP_TMPL3),

	.APUFCMDECFPUOP (APUFCMDECFPUOP_delay),
	.APUFCMDECLDSTXFERSIZE (APUFCMDECLDSTXFERSIZE_delay),
	.APUFCMDECLOAD (APUFCMDECLOAD_delay),
	.APUFCMDECNONAUTON (APUFCMDECNONAUTON_delay),
	.APUFCMDECSTORE (APUFCMDECSTORE_delay),
	.APUFCMDECUDI (APUFCMDECUDI_delay),
	.APUFCMDECUDIVALID (APUFCMDECUDIVALID_delay),
	.APUFCMENDIAN (APUFCMENDIAN_delay),
	.APUFCMFLUSH (APUFCMFLUSH_delay),
	.APUFCMINSTRUCTION (APUFCMINSTRUCTION_delay),
	.APUFCMINSTRVALID (APUFCMINSTRVALID_delay),
	.APUFCMLOADBYTEADDR (APUFCMLOADBYTEADDR_delay),
	.APUFCMLOADDATA (APUFCMLOADDATA_delay),
	.APUFCMLOADDVALID (APUFCMLOADDVALID_delay),
	.APUFCMMSRFE0 (APUFCMMSRFE0_delay),
	.APUFCMMSRFE1 (APUFCMMSRFE1_delay),
	.APUFCMNEXTINSTRREADY (APUFCMNEXTINSTRREADY_delay),
	.APUFCMOPERANDVALID (APUFCMOPERANDVALID_delay),
	.APUFCMRADATA (APUFCMRADATA_delay),
	.APUFCMRBDATA (APUFCMRBDATA_delay),
	.APUFCMWRITEBACKOK (APUFCMWRITEBACKOK_delay),
	.C440CPMCORESLEEPREQ (C440CPMCORESLEEPREQ_delay),
	.C440CPMDECIRPTREQ (C440CPMDECIRPTREQ_delay),
	.C440CPMFITIRPTREQ (C440CPMFITIRPTREQ_delay),
	.C440CPMMSRCE (C440CPMMSRCE_delay),
	.C440CPMMSREE (C440CPMMSREE_delay),
	.C440CPMTIMERRESETREQ (C440CPMTIMERRESETREQ_delay),
	.C440CPMWDIRPTREQ (C440CPMWDIRPTREQ_delay),
	.C440DBGSYSTEMCONTROL (C440DBGSYSTEMCONTROL_delay),
	.C440JTGTDO (C440JTGTDO_delay),
	.C440JTGTDOEN (C440JTGTDOEN_delay),
	.C440MACHINECHECK (C440MACHINECHECK_delay),
	.C440RSTCHIPRESETREQ (C440RSTCHIPRESETREQ_delay),
	.C440RSTCORERESETREQ (C440RSTCORERESETREQ_delay),
	.C440RSTSYSTEMRESETREQ (C440RSTSYSTEMRESETREQ_delay),
	.C440TRCBRANCHSTATUS (C440TRCBRANCHSTATUS_delay),
	.C440TRCCYCLE (C440TRCCYCLE_delay),
	.C440TRCEXECUTIONSTATUS (C440TRCEXECUTIONSTATUS_delay),
	.C440TRCTRACESTATUS (C440TRCTRACESTATUS_delay),
	.C440TRCTRIGGEREVENTOUT (C440TRCTRIGGEREVENTOUT_delay),
	.C440TRCTRIGGEREVENTTYPE (C440TRCTRIGGEREVENTTYPE_delay),
	.DMA0LLRSTENGINEACK (DMA0LLRSTENGINEACK_delay),
	.DMA0LLRXDSTRDYN (DMA0LLRXDSTRDYN_delay),
	.DMA0LLTXD (DMA0LLTXD_delay),
	.DMA0LLTXEOFN (DMA0LLTXEOFN_delay),
	.DMA0LLTXEOPN (DMA0LLTXEOPN_delay),
	.DMA0LLTXREM (DMA0LLTXREM_delay),
	.DMA0LLTXSOFN (DMA0LLTXSOFN_delay),
	.DMA0LLTXSOPN (DMA0LLTXSOPN_delay),
	.DMA0LLTXSRCRDYN (DMA0LLTXSRCRDYN_delay),
	.DMA0RXIRQ (DMA0RXIRQ_delay),
	.DMA0TXIRQ (DMA0TXIRQ_delay),
	.DMA1LLRSTENGINEACK (DMA1LLRSTENGINEACK_delay),
	.DMA1LLRXDSTRDYN (DMA1LLRXDSTRDYN_delay),
	.DMA1LLTXD (DMA1LLTXD_delay),
	.DMA1LLTXEOFN (DMA1LLTXEOFN_delay),
	.DMA1LLTXEOPN (DMA1LLTXEOPN_delay),
	.DMA1LLTXREM (DMA1LLTXREM_delay),
	.DMA1LLTXSOFN (DMA1LLTXSOFN_delay),
	.DMA1LLTXSOPN (DMA1LLTXSOPN_delay),
	.DMA1LLTXSRCRDYN (DMA1LLTXSRCRDYN_delay),
	.DMA1RXIRQ (DMA1RXIRQ_delay),
	.DMA1TXIRQ (DMA1TXIRQ_delay),
	.DMA2LLRSTENGINEACK (DMA2LLRSTENGINEACK_delay),
	.DMA2LLRXDSTRDYN (DMA2LLRXDSTRDYN_delay),
	.DMA2LLTXD (DMA2LLTXD_delay),
	.DMA2LLTXEOFN (DMA2LLTXEOFN_delay),
	.DMA2LLTXEOPN (DMA2LLTXEOPN_delay),
	.DMA2LLTXREM (DMA2LLTXREM_delay),
	.DMA2LLTXSOFN (DMA2LLTXSOFN_delay),
	.DMA2LLTXSOPN (DMA2LLTXSOPN_delay),
	.DMA2LLTXSRCRDYN (DMA2LLTXSRCRDYN_delay),
	.DMA2RXIRQ (DMA2RXIRQ_delay),
	.DMA2TXIRQ (DMA2TXIRQ_delay),
	.DMA3LLRSTENGINEACK (DMA3LLRSTENGINEACK_delay),
	.DMA3LLRXDSTRDYN (DMA3LLRXDSTRDYN_delay),
	.DMA3LLTXD (DMA3LLTXD_delay),
	.DMA3LLTXEOFN (DMA3LLTXEOFN_delay),
	.DMA3LLTXEOPN (DMA3LLTXEOPN_delay),
	.DMA3LLTXREM (DMA3LLTXREM_delay),
	.DMA3LLTXSOFN (DMA3LLTXSOFN_delay),
	.DMA3LLTXSOPN (DMA3LLTXSOPN_delay),
	.DMA3LLTXSRCRDYN (DMA3LLTXSRCRDYN_delay),
	.DMA3RXIRQ (DMA3RXIRQ_delay),
	.DMA3TXIRQ (DMA3TXIRQ_delay),
	.MIMCADDRESS (MIMCADDRESS_delay),
	.MIMCADDRESSVALID (MIMCADDRESSVALID_delay),
	.MIMCBANKCONFLICT (MIMCBANKCONFLICT_delay),
	.MIMCBYTEENABLE (MIMCBYTEENABLE_delay),
	.MIMCREADNOTWRITE (MIMCREADNOTWRITE_delay),
	.MIMCROWCONFLICT (MIMCROWCONFLICT_delay),
	.MIMCWRITEDATA (MIMCWRITEDATA_delay),
	.MIMCWRITEDATAVALID (MIMCWRITEDATAVALID_delay),
	.PPCCPMINTERCONNECTBUSY (PPCCPMINTERCONNECTBUSY_delay),
	.PPCDMDCRABUS (PPCDMDCRABUS_delay),
	.PPCDMDCRDBUSOUT (PPCDMDCRDBUSOUT_delay),
	.PPCDMDCRREAD (PPCDMDCRREAD_delay),
	.PPCDMDCRUABUS (PPCDMDCRUABUS_delay),
	.PPCDMDCRWRITE (PPCDMDCRWRITE_delay),
	.PPCDSDCRACK (PPCDSDCRACK_delay),
	.PPCDSDCRDBUSIN (PPCDSDCRDBUSIN_delay),
	.PPCDSDCRTIMEOUTWAIT (PPCDSDCRTIMEOUTWAIT_delay),
	.PPCEICINTERCONNECTIRQ (PPCEICINTERCONNECTIRQ_delay),
	.PPCMPLBABORT (PPCMPLBABORT_delay),
	.PPCMPLBABUS (PPCMPLBABUS_delay),
	.PPCMPLBBE (PPCMPLBBE_delay),
	.PPCMPLBBUSLOCK (PPCMPLBBUSLOCK_delay),
	.PPCMPLBLOCKERR (PPCMPLBLOCKERR_delay),
	.PPCMPLBPRIORITY (PPCMPLBPRIORITY_delay),
	.PPCMPLBRDBURST (PPCMPLBRDBURST_delay),
	.PPCMPLBREQUEST (PPCMPLBREQUEST_delay),
	.PPCMPLBRNW (PPCMPLBRNW_delay),
	.PPCMPLBSIZE (PPCMPLBSIZE_delay),
	.PPCMPLBTATTRIBUTE (PPCMPLBTATTRIBUTE_delay),
	.PPCMPLBTYPE (PPCMPLBTYPE_delay),
	.PPCMPLBUABUS (PPCMPLBUABUS_delay),
	.PPCMPLBWRBURST (PPCMPLBWRBURST_delay),
	.PPCMPLBWRDBUS (PPCMPLBWRDBUS_delay),
	.PPCS0PLBADDRACK (PPCS0PLBADDRACK_delay),
	.PPCS0PLBMBUSY (PPCS0PLBMBUSY_delay),
	.PPCS0PLBMIRQ (PPCS0PLBMIRQ_delay),
	.PPCS0PLBMRDERR (PPCS0PLBMRDERR_delay),
	.PPCS0PLBMWRERR (PPCS0PLBMWRERR_delay),
	.PPCS0PLBRDBTERM (PPCS0PLBRDBTERM_delay),
	.PPCS0PLBRDCOMP (PPCS0PLBRDCOMP_delay),
	.PPCS0PLBRDDACK (PPCS0PLBRDDACK_delay),
	.PPCS0PLBRDDBUS (PPCS0PLBRDDBUS_delay),
	.PPCS0PLBRDWDADDR (PPCS0PLBRDWDADDR_delay),
	.PPCS0PLBREARBITRATE (PPCS0PLBREARBITRATE_delay),
	.PPCS0PLBSSIZE (PPCS0PLBSSIZE_delay),
	.PPCS0PLBWAIT (PPCS0PLBWAIT_delay),
	.PPCS0PLBWRBTERM (PPCS0PLBWRBTERM_delay),
	.PPCS0PLBWRCOMP (PPCS0PLBWRCOMP_delay),
	.PPCS0PLBWRDACK (PPCS0PLBWRDACK_delay),
	.PPCS1PLBADDRACK (PPCS1PLBADDRACK_delay),
	.PPCS1PLBMBUSY (PPCS1PLBMBUSY_delay),
	.PPCS1PLBMIRQ (PPCS1PLBMIRQ_delay),
	.PPCS1PLBMRDERR (PPCS1PLBMRDERR_delay),
	.PPCS1PLBMWRERR (PPCS1PLBMWRERR_delay),
	.PPCS1PLBRDBTERM (PPCS1PLBRDBTERM_delay),
	.PPCS1PLBRDCOMP (PPCS1PLBRDCOMP_delay),
	.PPCS1PLBRDDACK (PPCS1PLBRDDACK_delay),
	.PPCS1PLBRDDBUS (PPCS1PLBRDDBUS_delay),
	.PPCS1PLBRDWDADDR (PPCS1PLBRDWDADDR_delay),
	.PPCS1PLBREARBITRATE (PPCS1PLBREARBITRATE_delay),
	.PPCS1PLBSSIZE (PPCS1PLBSSIZE_delay),
	.PPCS1PLBWAIT (PPCS1PLBWAIT_delay),
	.PPCS1PLBWRBTERM (PPCS1PLBWRBTERM_delay),
	.PPCS1PLBWRCOMP (PPCS1PLBWRCOMP_delay),
	.PPCS1PLBWRDACK (PPCS1PLBWRDACK_delay),

	.CPMC440CLK (CPMC440CLK_delay),
	.CPMC440CLKEN (CPMC440CLKEN_delay),
	.CPMC440CORECLOCKINACTIVE (CPMC440CORECLOCKINACTIVE_delay),
	.CPMC440TIMERCLOCK (CPMC440TIMERCLOCK_delay),
	.CPMDCRCLK (CPMDCRCLK_delay),
	.CPMDMA0LLCLK (CPMDMA0LLCLK_delay),
	.CPMDMA1LLCLK (CPMDMA1LLCLK_delay),
	.CPMDMA2LLCLK (CPMDMA2LLCLK_delay),
	.CPMDMA3LLCLK (CPMDMA3LLCLK_delay),
	.CPMFCMCLK (CPMFCMCLK_delay),
	.CPMINTERCONNECTCLK (CPMINTERCONNECTCLK_delay),
	.CPMINTERCONNECTCLKEN (CPMINTERCONNECTCLKEN_delay),
	.CPMINTERCONNECTCLKNTO1 (CPMINTERCONNECTCLKNTO1_delay),
	.CPMMCCLK (CPMMCCLK_delay),
	.CPMPPCMPLBCLK (CPMPPCMPLBCLK_delay),
	.CPMPPCS0PLBCLK (CPMPPCS0PLBCLK_delay),
	.CPMPPCS1PLBCLK (CPMPPCS1PLBCLK_delay),
	.DBGC440DEBUGHALT (DBGC440DEBUGHALT_delay),
	.DBGC440SYSTEMSTATUS (DBGC440SYSTEMSTATUS_delay),
	.DBGC440UNCONDDEBUGEVENT (DBGC440UNCONDDEBUGEVENT_delay),
	.DCRPPCDMACK (DCRPPCDMACK_delay),
	.DCRPPCDMDBUSIN (DCRPPCDMDBUSIN_delay),
	.DCRPPCDMTIMEOUTWAIT (DCRPPCDMTIMEOUTWAIT_delay),
	.DCRPPCDSABUS (DCRPPCDSABUS_delay),
	.DCRPPCDSDBUSOUT (DCRPPCDSDBUSOUT_delay),
	.DCRPPCDSREAD (DCRPPCDSREAD_delay),
	.DCRPPCDSWRITE (DCRPPCDSWRITE_delay),
	.EICC440CRITIRQ (EICC440CRITIRQ_delay),
	.EICC440EXTIRQ (EICC440EXTIRQ_delay),
	.FCMAPUCONFIRMINSTR (FCMAPUCONFIRMINSTR_delay),
	.FCMAPUCR (FCMAPUCR_delay),
	.FCMAPUDONE (FCMAPUDONE_delay),
	.FCMAPUEXCEPTION (FCMAPUEXCEPTION_delay),
	.FCMAPUFPSCRFEX (FCMAPUFPSCRFEX_delay),
	.FCMAPURESULT (FCMAPURESULT_delay),
	.FCMAPURESULTVALID (FCMAPURESULTVALID_delay),
	.FCMAPUSLEEPNOTREADY (FCMAPUSLEEPNOTREADY_delay),
	.FCMAPUSTOREDATA (FCMAPUSTOREDATA_delay),
	.JTGC440TCK (JTGC440TCK_delay),
	.JTGC440TDI (JTGC440TDI_delay),
	.JTGC440TMS (JTGC440TMS_delay),
	.JTGC440TRSTNEG (JTGC440TRSTNEG_delay),
	.LLDMA0RSTENGINEREQ (LLDMA0RSTENGINEREQ_delay),
	.LLDMA0RXD (LLDMA0RXD_delay),
	.LLDMA0RXEOFN (LLDMA0RXEOFN_delay),
	.LLDMA0RXEOPN (LLDMA0RXEOPN_delay),
	.LLDMA0RXREM (LLDMA0RXREM_delay),
	.LLDMA0RXSOFN (LLDMA0RXSOFN_delay),
	.LLDMA0RXSOPN (LLDMA0RXSOPN_delay),
	.LLDMA0RXSRCRDYN (LLDMA0RXSRCRDYN_delay),
	.LLDMA0TXDSTRDYN (LLDMA0TXDSTRDYN_delay),
	.LLDMA1RSTENGINEREQ (LLDMA1RSTENGINEREQ_delay),
	.LLDMA1RXD (LLDMA1RXD_delay),
	.LLDMA1RXEOFN (LLDMA1RXEOFN_delay),
	.LLDMA1RXEOPN (LLDMA1RXEOPN_delay),
	.LLDMA1RXREM (LLDMA1RXREM_delay),
	.LLDMA1RXSOFN (LLDMA1RXSOFN_delay),
	.LLDMA1RXSOPN (LLDMA1RXSOPN_delay),
	.LLDMA1RXSRCRDYN (LLDMA1RXSRCRDYN_delay),
	.LLDMA1TXDSTRDYN (LLDMA1TXDSTRDYN_delay),
	.LLDMA2RSTENGINEREQ (LLDMA2RSTENGINEREQ_delay),
	.LLDMA2RXD (LLDMA2RXD_delay),
	.LLDMA2RXEOFN (LLDMA2RXEOFN_delay),
	.LLDMA2RXEOPN (LLDMA2RXEOPN_delay),
	.LLDMA2RXREM (LLDMA2RXREM_delay),
	.LLDMA2RXSOFN (LLDMA2RXSOFN_delay),
	.LLDMA2RXSOPN (LLDMA2RXSOPN_delay),
	.LLDMA2RXSRCRDYN (LLDMA2RXSRCRDYN_delay),
	.LLDMA2TXDSTRDYN (LLDMA2TXDSTRDYN_delay),
	.LLDMA3RSTENGINEREQ (LLDMA3RSTENGINEREQ_delay),
	.LLDMA3RXD (LLDMA3RXD_delay),
	.LLDMA3RXEOFN (LLDMA3RXEOFN_delay),
	.LLDMA3RXEOPN (LLDMA3RXEOPN_delay),
	.LLDMA3RXREM (LLDMA3RXREM_delay),
	.LLDMA3RXSOFN (LLDMA3RXSOFN_delay),
	.LLDMA3RXSOPN (LLDMA3RXSOPN_delay),
	.LLDMA3RXSRCRDYN (LLDMA3RXSRCRDYN_delay),
	.LLDMA3TXDSTRDYN (LLDMA3TXDSTRDYN_delay),
	.MCMIADDRREADYTOACCEPT (MCMIADDRREADYTOACCEPT_delay),
	.MCMIREADDATA (MCMIREADDATA_delay),
	.MCMIREADDATAERR (MCMIREADDATAERR_delay),
	.MCMIREADDATAVALID (MCMIREADDATAVALID_delay),
	.PLBPPCMADDRACK (PLBPPCMADDRACK_delay),
	.PLBPPCMMBUSY (PLBPPCMMBUSY_delay),
	.PLBPPCMMIRQ (PLBPPCMMIRQ_delay),
	.PLBPPCMMRDERR (PLBPPCMMRDERR_delay),
	.PLBPPCMMWRERR (PLBPPCMMWRERR_delay),
	.PLBPPCMRDBTERM (PLBPPCMRDBTERM_delay),
	.PLBPPCMRDDACK (PLBPPCMRDDACK_delay),
	.PLBPPCMRDDBUS (PLBPPCMRDDBUS_delay),
	.PLBPPCMRDPENDPRI (PLBPPCMRDPENDPRI_delay),
	.PLBPPCMRDPENDREQ (PLBPPCMRDPENDREQ_delay),
	.PLBPPCMRDWDADDR (PLBPPCMRDWDADDR_delay),
	.PLBPPCMREARBITRATE (PLBPPCMREARBITRATE_delay),
	.PLBPPCMREQPRI (PLBPPCMREQPRI_delay),
	.PLBPPCMSSIZE (PLBPPCMSSIZE_delay),
	.PLBPPCMTIMEOUT (PLBPPCMTIMEOUT_delay),
	.PLBPPCMWRBTERM (PLBPPCMWRBTERM_delay),
	.PLBPPCMWRDACK (PLBPPCMWRDACK_delay),
	.PLBPPCMWRPENDPRI (PLBPPCMWRPENDPRI_delay),
	.PLBPPCMWRPENDREQ (PLBPPCMWRPENDREQ_delay),
	.PLBPPCS0ABORT (PLBPPCS0ABORT_delay),
	.PLBPPCS0ABUS (PLBPPCS0ABUS_delay),
	.PLBPPCS0BE (PLBPPCS0BE_delay),
	.PLBPPCS0BUSLOCK (PLBPPCS0BUSLOCK_delay),
	.PLBPPCS0LOCKERR (PLBPPCS0LOCKERR_delay),
	.PLBPPCS0MASTERID (PLBPPCS0MASTERID_delay),
	.PLBPPCS0MSIZE (PLBPPCS0MSIZE_delay),
	.PLBPPCS0PAVALID (PLBPPCS0PAVALID_delay),
	.PLBPPCS0RDBURST (PLBPPCS0RDBURST_delay),
	.PLBPPCS0RDPENDPRI (PLBPPCS0RDPENDPRI_delay),
	.PLBPPCS0RDPENDREQ (PLBPPCS0RDPENDREQ_delay),
	.PLBPPCS0RDPRIM (PLBPPCS0RDPRIM_delay),
	.PLBPPCS0REQPRI (PLBPPCS0REQPRI_delay),
	.PLBPPCS0RNW (PLBPPCS0RNW_delay),
	.PLBPPCS0SAVALID (PLBPPCS0SAVALID_delay),
	.PLBPPCS0SIZE (PLBPPCS0SIZE_delay),
	.PLBPPCS0TATTRIBUTE (PLBPPCS0TATTRIBUTE_delay),
	.PLBPPCS0TYPE (PLBPPCS0TYPE_delay),
	.PLBPPCS0UABUS (PLBPPCS0UABUS_delay),
	.PLBPPCS0WRBURST (PLBPPCS0WRBURST_delay),
	.PLBPPCS0WRDBUS (PLBPPCS0WRDBUS_delay),
	.PLBPPCS0WRPENDPRI (PLBPPCS0WRPENDPRI_delay),
	.PLBPPCS0WRPENDREQ (PLBPPCS0WRPENDREQ_delay),
	.PLBPPCS0WRPRIM (PLBPPCS0WRPRIM_delay),
	.PLBPPCS1ABORT (PLBPPCS1ABORT_delay),
	.PLBPPCS1ABUS (PLBPPCS1ABUS_delay),
	.PLBPPCS1BE (PLBPPCS1BE_delay),
	.PLBPPCS1BUSLOCK (PLBPPCS1BUSLOCK_delay),
	.PLBPPCS1LOCKERR (PLBPPCS1LOCKERR_delay),
	.PLBPPCS1MASTERID (PLBPPCS1MASTERID_delay),
	.PLBPPCS1MSIZE (PLBPPCS1MSIZE_delay),
	.PLBPPCS1PAVALID (PLBPPCS1PAVALID_delay),
	.PLBPPCS1RDBURST (PLBPPCS1RDBURST_delay),
	.PLBPPCS1RDPENDPRI (PLBPPCS1RDPENDPRI_delay),
	.PLBPPCS1RDPENDREQ (PLBPPCS1RDPENDREQ_delay),
	.PLBPPCS1RDPRIM (PLBPPCS1RDPRIM_delay),
	.PLBPPCS1REQPRI (PLBPPCS1REQPRI_delay),
	.PLBPPCS1RNW (PLBPPCS1RNW_delay),
	.PLBPPCS1SAVALID (PLBPPCS1SAVALID_delay),
	.PLBPPCS1SIZE (PLBPPCS1SIZE_delay),
	.PLBPPCS1TATTRIBUTE (PLBPPCS1TATTRIBUTE_delay),
	.PLBPPCS1TYPE (PLBPPCS1TYPE_delay),
	.PLBPPCS1UABUS (PLBPPCS1UABUS_delay),
	.PLBPPCS1WRBURST (PLBPPCS1WRBURST_delay),
	.PLBPPCS1WRDBUS (PLBPPCS1WRDBUS_delay),
	.PLBPPCS1WRPENDPRI (PLBPPCS1WRPENDPRI_delay),
	.PLBPPCS1WRPENDREQ (PLBPPCS1WRPENDREQ_delay),
	.PLBPPCS1WRPRIM (PLBPPCS1WRPRIM_delay),
	.RSTC440RESETCHIP (RSTC440RESETCHIP_delay),
	.RSTC440RESETCORE (RSTC440RESETCORE_delay),
	.RSTC440RESETSYSTEM (RSTC440RESETSYSTEM_delay),
	.TIEC440DCURDLDCACHEPLBPRIO (TIEC440DCURDLDCACHEPLBPRIO_delay),
	.TIEC440DCURDNONCACHEPLBPRIO (TIEC440DCURDNONCACHEPLBPRIO_delay),
	.TIEC440DCURDTOUCHPLBPRIO (TIEC440DCURDTOUCHPLBPRIO_delay),
	.TIEC440DCURDURGENTPLBPRIO (TIEC440DCURDURGENTPLBPRIO_delay),
	.TIEC440DCUWRFLUSHPLBPRIO (TIEC440DCUWRFLUSHPLBPRIO_delay),
	.TIEC440DCUWRSTOREPLBPRIO (TIEC440DCUWRSTOREPLBPRIO_delay),
	.TIEC440DCUWRURGENTPLBPRIO (TIEC440DCUWRURGENTPLBPRIO_delay),
	.TIEC440ENDIANRESET (TIEC440ENDIANRESET_delay),
	.TIEC440ERPNRESET (TIEC440ERPNRESET_delay),
	.TIEC440ICURDFETCHPLBPRIO (TIEC440ICURDFETCHPLBPRIO_delay),
	.TIEC440ICURDSPECPLBPRIO (TIEC440ICURDSPECPLBPRIO_delay),
	.TIEC440ICURDTOUCHPLBPRIO (TIEC440ICURDTOUCHPLBPRIO_delay),
	.TIEC440PIR (TIEC440PIR_delay),
	.TIEC440PVR (TIEC440PVR_delay),
	.TIEC440USERRESET (TIEC440USERRESET_delay),
	.TIEDCRBASEADDR (TIEDCRBASEADDR_delay),
	.TRCC440TRACEDISABLE (TRCC440TRACEDISABLE_delay),
	.TRCC440TRIGGEREVENTIN (TRCC440TRIGGEREVENTIN_delay),
	.GSR (GSR)
);

specify
	$period (posedge CPMC440TIMERCLOCK, 0:0:0);
	$period (posedge CPMDCRCLK, 0:0:0);
	$period (posedge CPMFCMCLK, 0:0:0);
	$period (posedge CPMINTERCONNECTCLK, 0:0:0);
	$period (posedge CPMMCCLK, 0:0:0);
	$period (posedge CPMPPCMPLBCLK, 0:0:0);
	$period (posedge CPMPPCS0PLBCLK, 0:0:0);
	$period (posedge CPMPPCS1PLBCLK, 0:0:0);
	$setuphold (posedge CPMC440CLK, negedge DBGC440DEBUGHALT, 0:0:0, 0:0:0, notifier,,,CPMC440CLK_delay,DBGC440DEBUGHALT_delay);
	$setuphold (posedge CPMC440CLK, negedge DBGC440UNCONDDEBUGEVENT, 0:0:0, 0:0:0, notifier,,,CPMC440CLK_delay,DBGC440UNCONDDEBUGEVENT_delay);
	$setuphold (posedge CPMC440CLK, negedge TRCC440TRACEDISABLE, 0:0:0, 0:0:0, notifier,,,CPMC440CLK_delay,TRCC440TRACEDISABLE_delay);
	$setuphold (posedge CPMC440CLK, negedge TRCC440TRIGGEREVENTIN, 0:0:0, 0:0:0, notifier,,,CPMC440CLK_delay,TRCC440TRIGGEREVENTIN_delay);
	$setuphold (posedge CPMC440CLK, posedge DBGC440DEBUGHALT, 0:0:0, 0:0:0, notifier,,,CPMC440CLK_delay,DBGC440DEBUGHALT_delay);
	$setuphold (posedge CPMC440CLK, posedge DBGC440UNCONDDEBUGEVENT, 0:0:0, 0:0:0, notifier,,,CPMC440CLK_delay,DBGC440UNCONDDEBUGEVENT_delay);
	$setuphold (posedge CPMC440CLK, posedge TRCC440TRACEDISABLE, 0:0:0, 0:0:0, notifier,,,CPMC440CLK_delay,TRCC440TRACEDISABLE_delay);
	$setuphold (posedge CPMC440CLK, posedge TRCC440TRIGGEREVENTIN, 0:0:0, 0:0:0, notifier,,,CPMC440CLK_delay,TRCC440TRIGGEREVENTIN_delay);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMACK, 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMACK_delay);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[0], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[0]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[10], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[10]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[11], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[11]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[12], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[12]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[13], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[13]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[14], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[14]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[15], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[15]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[16], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[16]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[17], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[17]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[18], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[18]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[19], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[19]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[1], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[1]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[20], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[20]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[21], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[21]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[22], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[22]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[23], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[23]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[24], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[24]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[25], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[25]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[26], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[26]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[27], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[27]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[28], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[28]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[29], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[29]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[2], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[2]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[30], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[30]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[31], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[31]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[3], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[3]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[4], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[4]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[5], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[5]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[6], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[6]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[7], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[7]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[8], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[8]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMDBUSIN[9], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[9]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDMTIMEOUTWAIT, 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMTIMEOUTWAIT_delay);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSABUS[0], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[0]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSABUS[1], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[1]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSABUS[2], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[2]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSABUS[3], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[3]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSABUS[4], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[4]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSABUS[5], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[5]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSABUS[6], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[6]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSABUS[7], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[7]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSABUS[8], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[8]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSABUS[9], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[9]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[0], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[0]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[10], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[10]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[11], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[11]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[12], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[12]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[13], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[13]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[14], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[14]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[15], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[15]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[16], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[16]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[17], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[17]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[18], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[18]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[19], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[19]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[1], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[1]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[20], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[20]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[21], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[21]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[22], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[22]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[23], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[23]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[24], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[24]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[25], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[25]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[26], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[26]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[27], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[27]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[28], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[28]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[29], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[29]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[2], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[2]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[30], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[30]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[31], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[31]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[3], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[3]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[4], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[4]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[5], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[5]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[6], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[6]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[7], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[7]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[8], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[8]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSDBUSOUT[9], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[9]);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSREAD, 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSREAD_delay);
	$setuphold (posedge CPMDCRCLK, negedge DCRPPCDSWRITE, 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSWRITE_delay);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMACK, 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMACK_delay);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[0], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[0]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[10], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[10]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[11], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[11]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[12], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[12]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[13], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[13]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[14], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[14]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[15], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[15]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[16], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[16]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[17], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[17]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[18], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[18]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[19], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[19]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[1], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[1]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[20], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[20]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[21], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[21]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[22], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[22]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[23], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[23]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[24], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[24]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[25], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[25]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[26], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[26]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[27], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[27]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[28], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[28]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[29], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[29]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[2], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[2]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[30], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[30]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[31], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[31]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[3], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[3]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[4], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[4]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[5], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[5]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[6], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[6]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[7], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[7]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[8], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[8]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMDBUSIN[9], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMDBUSIN_delay[9]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDMTIMEOUTWAIT, 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDMTIMEOUTWAIT_delay);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSABUS[0], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[0]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSABUS[1], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[1]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSABUS[2], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[2]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSABUS[3], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[3]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSABUS[4], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[4]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSABUS[5], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[5]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSABUS[6], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[6]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSABUS[7], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[7]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSABUS[8], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[8]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSABUS[9], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSABUS_delay[9]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[0], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[0]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[10], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[10]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[11], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[11]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[12], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[12]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[13], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[13]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[14], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[14]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[15], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[15]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[16], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[16]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[17], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[17]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[18], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[18]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[19], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[19]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[1], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[1]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[20], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[20]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[21], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[21]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[22], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[22]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[23], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[23]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[24], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[24]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[25], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[25]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[26], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[26]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[27], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[27]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[28], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[28]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[29], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[29]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[2], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[2]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[30], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[30]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[31], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[31]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[3], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[3]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[4], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[4]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[5], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[5]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[6], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[6]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[7], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[7]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[8], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[8]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSDBUSOUT[9], 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSDBUSOUT_delay[9]);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSREAD, 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSREAD_delay);
	$setuphold (posedge CPMDCRCLK, posedge DCRPPCDSWRITE, 0:0:0, 0:0:0, notifier,,,CPMDCRCLK_delay,DCRPPCDSWRITE_delay);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RSTENGINEREQ, 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RSTENGINEREQ_delay);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[0], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[0]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[10], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[10]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[11], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[11]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[12], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[12]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[13], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[13]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[14], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[14]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[15], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[15]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[16], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[16]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[17], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[17]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[18], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[18]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[19], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[19]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[1], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[1]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[20], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[20]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[21], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[21]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[22], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[22]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[23], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[23]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[24], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[24]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[25], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[25]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[26], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[26]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[27], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[27]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[28], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[28]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[29], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[29]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[2], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[2]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[30], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[30]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[31], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[31]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[3], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[3]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[4], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[4]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[5], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[5]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[6], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[6]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[7], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[7]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[8], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[8]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXD[9], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[9]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXEOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXEOFN_delay);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXEOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXEOPN_delay);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXREM[0], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXREM_delay[0]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXREM[1], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXREM_delay[1]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXREM[2], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXREM_delay[2]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXREM[3], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXREM_delay[3]);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXSOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXSOFN_delay);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXSOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXSOPN_delay);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0RXSRCRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXSRCRDYN_delay);
	$setuphold (posedge CPMDMA0LLCLK, negedge LLDMA0TXDSTRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0TXDSTRDYN_delay);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RSTENGINEREQ, 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RSTENGINEREQ_delay);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[0], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[0]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[10], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[10]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[11], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[11]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[12], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[12]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[13], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[13]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[14], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[14]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[15], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[15]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[16], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[16]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[17], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[17]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[18], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[18]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[19], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[19]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[1], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[1]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[20], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[20]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[21], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[21]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[22], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[22]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[23], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[23]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[24], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[24]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[25], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[25]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[26], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[26]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[27], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[27]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[28], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[28]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[29], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[29]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[2], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[2]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[30], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[30]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[31], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[31]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[3], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[3]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[4], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[4]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[5], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[5]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[6], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[6]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[7], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[7]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[8], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[8]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXD[9], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXD_delay[9]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXEOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXEOFN_delay);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXEOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXEOPN_delay);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXREM[0], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXREM_delay[0]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXREM[1], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXREM_delay[1]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXREM[2], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXREM_delay[2]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXREM[3], 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXREM_delay[3]);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXSOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXSOFN_delay);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXSOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXSOPN_delay);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0RXSRCRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0RXSRCRDYN_delay);
	$setuphold (posedge CPMDMA0LLCLK, posedge LLDMA0TXDSTRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA0LLCLK_delay,LLDMA0TXDSTRDYN_delay);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RSTENGINEREQ, 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RSTENGINEREQ_delay);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[0], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[0]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[10], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[10]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[11], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[11]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[12], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[12]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[13], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[13]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[14], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[14]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[15], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[15]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[16], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[16]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[17], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[17]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[18], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[18]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[19], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[19]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[1], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[1]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[20], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[20]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[21], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[21]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[22], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[22]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[23], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[23]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[24], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[24]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[25], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[25]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[26], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[26]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[27], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[27]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[28], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[28]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[29], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[29]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[2], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[2]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[30], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[30]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[31], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[31]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[3], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[3]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[4], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[4]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[5], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[5]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[6], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[6]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[7], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[7]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[8], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[8]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXD[9], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[9]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXEOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXEOFN_delay);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXEOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXEOPN_delay);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXREM[0], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXREM_delay[0]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXREM[1], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXREM_delay[1]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXREM[2], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXREM_delay[2]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXREM[3], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXREM_delay[3]);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXSOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXSOFN_delay);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXSOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXSOPN_delay);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1RXSRCRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXSRCRDYN_delay);
	$setuphold (posedge CPMDMA1LLCLK, negedge LLDMA1TXDSTRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1TXDSTRDYN_delay);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RSTENGINEREQ, 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RSTENGINEREQ_delay);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[0], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[0]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[10], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[10]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[11], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[11]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[12], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[12]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[13], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[13]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[14], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[14]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[15], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[15]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[16], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[16]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[17], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[17]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[18], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[18]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[19], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[19]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[1], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[1]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[20], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[20]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[21], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[21]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[22], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[22]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[23], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[23]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[24], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[24]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[25], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[25]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[26], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[26]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[27], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[27]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[28], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[28]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[29], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[29]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[2], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[2]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[30], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[30]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[31], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[31]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[3], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[3]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[4], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[4]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[5], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[5]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[6], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[6]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[7], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[7]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[8], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[8]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXD[9], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXD_delay[9]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXEOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXEOFN_delay);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXEOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXEOPN_delay);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXREM[0], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXREM_delay[0]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXREM[1], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXREM_delay[1]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXREM[2], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXREM_delay[2]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXREM[3], 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXREM_delay[3]);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXSOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXSOFN_delay);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXSOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXSOPN_delay);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1RXSRCRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1RXSRCRDYN_delay);
	$setuphold (posedge CPMDMA1LLCLK, posedge LLDMA1TXDSTRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA1LLCLK_delay,LLDMA1TXDSTRDYN_delay);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RSTENGINEREQ, 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RSTENGINEREQ_delay);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[0], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[0]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[10], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[10]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[11], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[11]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[12], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[12]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[13], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[13]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[14], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[14]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[15], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[15]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[16], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[16]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[17], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[17]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[18], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[18]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[19], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[19]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[1], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[1]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[20], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[20]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[21], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[21]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[22], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[22]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[23], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[23]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[24], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[24]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[25], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[25]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[26], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[26]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[27], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[27]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[28], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[28]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[29], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[29]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[2], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[2]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[30], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[30]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[31], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[31]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[3], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[3]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[4], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[4]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[5], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[5]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[6], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[6]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[7], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[7]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[8], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[8]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXD[9], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[9]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXEOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXEOFN_delay);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXEOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXEOPN_delay);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXREM[0], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXREM_delay[0]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXREM[1], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXREM_delay[1]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXREM[2], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXREM_delay[2]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXREM[3], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXREM_delay[3]);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXSOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXSOFN_delay);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXSOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXSOPN_delay);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2RXSRCRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXSRCRDYN_delay);
	$setuphold (posedge CPMDMA2LLCLK, negedge LLDMA2TXDSTRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2TXDSTRDYN_delay);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RSTENGINEREQ, 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RSTENGINEREQ_delay);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[0], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[0]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[10], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[10]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[11], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[11]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[12], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[12]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[13], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[13]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[14], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[14]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[15], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[15]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[16], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[16]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[17], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[17]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[18], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[18]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[19], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[19]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[1], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[1]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[20], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[20]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[21], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[21]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[22], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[22]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[23], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[23]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[24], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[24]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[25], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[25]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[26], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[26]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[27], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[27]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[28], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[28]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[29], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[29]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[2], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[2]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[30], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[30]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[31], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[31]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[3], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[3]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[4], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[4]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[5], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[5]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[6], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[6]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[7], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[7]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[8], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[8]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXD[9], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXD_delay[9]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXEOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXEOFN_delay);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXEOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXEOPN_delay);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXREM[0], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXREM_delay[0]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXREM[1], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXREM_delay[1]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXREM[2], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXREM_delay[2]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXREM[3], 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXREM_delay[3]);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXSOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXSOFN_delay);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXSOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXSOPN_delay);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2RXSRCRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2RXSRCRDYN_delay);
	$setuphold (posedge CPMDMA2LLCLK, posedge LLDMA2TXDSTRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA2LLCLK_delay,LLDMA2TXDSTRDYN_delay);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RSTENGINEREQ, 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RSTENGINEREQ_delay);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[0], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[0]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[10], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[10]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[11], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[11]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[12], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[12]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[13], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[13]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[14], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[14]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[15], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[15]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[16], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[16]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[17], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[17]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[18], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[18]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[19], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[19]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[1], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[1]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[20], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[20]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[21], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[21]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[22], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[22]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[23], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[23]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[24], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[24]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[25], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[25]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[26], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[26]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[27], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[27]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[28], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[28]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[29], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[29]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[2], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[2]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[30], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[30]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[31], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[31]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[3], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[3]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[4], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[4]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[5], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[5]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[6], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[6]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[7], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[7]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[8], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[8]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXD[9], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[9]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXEOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXEOFN_delay);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXEOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXEOPN_delay);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXREM[0], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXREM_delay[0]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXREM[1], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXREM_delay[1]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXREM[2], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXREM_delay[2]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXREM[3], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXREM_delay[3]);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXSOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXSOFN_delay);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXSOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXSOPN_delay);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3RXSRCRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXSRCRDYN_delay);
	$setuphold (posedge CPMDMA3LLCLK, negedge LLDMA3TXDSTRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3TXDSTRDYN_delay);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RSTENGINEREQ, 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RSTENGINEREQ_delay);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[0], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[0]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[10], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[10]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[11], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[11]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[12], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[12]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[13], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[13]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[14], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[14]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[15], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[15]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[16], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[16]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[17], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[17]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[18], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[18]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[19], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[19]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[1], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[1]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[20], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[20]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[21], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[21]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[22], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[22]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[23], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[23]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[24], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[24]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[25], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[25]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[26], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[26]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[27], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[27]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[28], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[28]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[29], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[29]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[2], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[2]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[30], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[30]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[31], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[31]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[3], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[3]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[4], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[4]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[5], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[5]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[6], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[6]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[7], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[7]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[8], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[8]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXD[9], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXD_delay[9]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXEOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXEOFN_delay);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXEOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXEOPN_delay);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXREM[0], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXREM_delay[0]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXREM[1], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXREM_delay[1]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXREM[2], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXREM_delay[2]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXREM[3], 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXREM_delay[3]);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXSOFN, 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXSOFN_delay);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXSOPN, 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXSOPN_delay);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3RXSRCRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3RXSRCRDYN_delay);
	$setuphold (posedge CPMDMA3LLCLK, posedge LLDMA3TXDSTRDYN, 0:0:0, 0:0:0, notifier,,,CPMDMA3LLCLK_delay,LLDMA3TXDSTRDYN_delay);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUCONFIRMINSTR, 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUCONFIRMINSTR_delay);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUCR[0], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUCR_delay[0]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUCR[1], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUCR_delay[1]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUCR[2], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUCR_delay[2]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUCR[3], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUCR_delay[3]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUDONE, 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUDONE_delay);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUEXCEPTION, 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUEXCEPTION_delay);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUFPSCRFEX, 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUFPSCRFEX_delay);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULTVALID, 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULTVALID_delay);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[0], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[0]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[10], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[10]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[11], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[11]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[12], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[12]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[13], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[13]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[14], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[14]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[15], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[15]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[16], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[16]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[17], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[17]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[18], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[18]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[19], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[19]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[1], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[1]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[20], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[20]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[21], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[21]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[22], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[22]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[23], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[23]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[24], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[24]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[25], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[25]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[26], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[26]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[27], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[27]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[28], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[28]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[29], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[29]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[2], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[2]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[30], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[30]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[31], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[31]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[3], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[3]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[4], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[4]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[5], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[5]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[6], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[6]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[7], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[7]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[8], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[8]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPURESULT[9], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[9]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSLEEPNOTREADY, 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSLEEPNOTREADY_delay);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[0], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[0]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[100], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[100]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[101], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[101]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[102], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[102]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[103], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[103]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[104], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[104]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[105], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[105]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[106], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[106]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[107], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[107]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[108], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[108]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[109], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[109]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[10], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[10]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[110], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[110]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[111], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[111]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[112], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[112]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[113], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[113]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[114], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[114]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[115], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[115]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[116], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[116]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[117], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[117]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[118], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[118]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[119], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[119]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[11], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[11]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[120], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[120]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[121], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[121]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[122], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[122]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[123], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[123]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[124], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[124]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[125], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[125]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[126], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[126]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[127], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[127]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[12], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[12]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[13], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[13]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[14], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[14]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[15], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[15]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[16], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[16]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[17], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[17]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[18], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[18]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[19], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[19]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[1], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[1]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[20], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[20]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[21], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[21]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[22], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[22]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[23], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[23]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[24], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[24]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[25], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[25]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[26], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[26]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[27], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[27]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[28], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[28]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[29], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[29]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[2], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[2]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[30], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[30]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[31], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[31]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[32], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[32]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[33], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[33]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[34], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[34]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[35], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[35]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[36], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[36]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[37], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[37]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[38], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[38]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[39], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[39]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[3], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[3]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[40], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[40]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[41], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[41]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[42], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[42]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[43], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[43]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[44], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[44]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[45], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[45]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[46], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[46]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[47], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[47]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[48], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[48]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[49], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[49]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[4], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[4]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[50], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[50]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[51], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[51]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[52], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[52]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[53], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[53]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[54], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[54]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[55], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[55]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[56], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[56]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[57], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[57]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[58], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[58]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[59], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[59]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[5], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[5]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[60], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[60]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[61], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[61]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[62], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[62]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[63], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[63]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[64], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[64]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[65], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[65]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[66], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[66]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[67], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[67]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[68], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[68]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[69], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[69]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[6], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[6]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[70], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[70]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[71], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[71]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[72], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[72]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[73], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[73]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[74], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[74]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[75], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[75]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[76], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[76]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[77], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[77]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[78], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[78]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[79], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[79]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[7], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[7]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[80], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[80]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[81], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[81]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[82], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[82]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[83], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[83]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[84], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[84]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[85], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[85]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[86], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[86]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[87], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[87]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[88], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[88]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[89], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[89]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[8], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[8]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[90], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[90]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[91], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[91]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[92], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[92]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[93], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[93]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[94], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[94]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[95], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[95]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[96], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[96]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[97], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[97]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[98], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[98]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[99], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[99]);
	$setuphold (posedge CPMFCMCLK, negedge FCMAPUSTOREDATA[9], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[9]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUCONFIRMINSTR, 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUCONFIRMINSTR_delay);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUCR[0], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUCR_delay[0]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUCR[1], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUCR_delay[1]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUCR[2], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUCR_delay[2]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUCR[3], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUCR_delay[3]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUDONE, 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUDONE_delay);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUEXCEPTION, 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUEXCEPTION_delay);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUFPSCRFEX, 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUFPSCRFEX_delay);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULTVALID, 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULTVALID_delay);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[0], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[0]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[10], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[10]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[11], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[11]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[12], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[12]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[13], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[13]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[14], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[14]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[15], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[15]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[16], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[16]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[17], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[17]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[18], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[18]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[19], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[19]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[1], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[1]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[20], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[20]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[21], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[21]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[22], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[22]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[23], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[23]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[24], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[24]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[25], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[25]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[26], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[26]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[27], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[27]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[28], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[28]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[29], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[29]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[2], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[2]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[30], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[30]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[31], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[31]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[3], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[3]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[4], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[4]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[5], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[5]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[6], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[6]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[7], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[7]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[8], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[8]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPURESULT[9], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPURESULT_delay[9]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSLEEPNOTREADY, 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSLEEPNOTREADY_delay);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[0], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[0]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[100], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[100]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[101], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[101]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[102], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[102]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[103], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[103]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[104], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[104]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[105], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[105]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[106], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[106]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[107], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[107]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[108], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[108]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[109], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[109]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[10], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[10]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[110], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[110]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[111], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[111]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[112], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[112]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[113], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[113]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[114], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[114]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[115], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[115]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[116], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[116]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[117], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[117]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[118], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[118]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[119], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[119]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[11], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[11]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[120], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[120]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[121], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[121]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[122], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[122]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[123], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[123]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[124], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[124]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[125], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[125]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[126], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[126]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[127], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[127]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[12], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[12]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[13], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[13]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[14], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[14]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[15], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[15]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[16], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[16]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[17], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[17]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[18], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[18]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[19], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[19]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[1], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[1]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[20], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[20]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[21], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[21]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[22], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[22]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[23], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[23]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[24], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[24]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[25], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[25]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[26], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[26]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[27], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[27]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[28], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[28]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[29], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[29]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[2], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[2]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[30], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[30]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[31], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[31]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[32], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[32]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[33], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[33]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[34], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[34]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[35], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[35]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[36], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[36]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[37], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[37]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[38], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[38]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[39], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[39]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[3], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[3]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[40], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[40]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[41], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[41]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[42], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[42]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[43], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[43]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[44], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[44]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[45], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[45]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[46], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[46]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[47], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[47]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[48], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[48]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[49], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[49]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[4], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[4]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[50], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[50]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[51], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[51]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[52], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[52]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[53], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[53]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[54], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[54]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[55], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[55]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[56], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[56]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[57], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[57]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[58], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[58]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[59], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[59]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[5], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[5]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[60], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[60]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[61], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[61]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[62], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[62]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[63], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[63]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[64], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[64]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[65], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[65]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[66], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[66]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[67], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[67]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[68], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[68]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[69], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[69]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[6], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[6]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[70], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[70]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[71], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[71]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[72], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[72]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[73], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[73]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[74], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[74]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[75], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[75]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[76], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[76]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[77], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[77]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[78], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[78]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[79], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[79]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[7], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[7]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[80], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[80]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[81], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[81]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[82], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[82]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[83], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[83]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[84], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[84]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[85], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[85]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[86], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[86]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[87], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[87]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[88], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[88]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[89], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[89]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[8], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[8]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[90], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[90]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[91], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[91]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[92], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[92]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[93], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[93]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[94], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[94]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[95], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[95]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[96], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[96]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[97], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[97]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[98], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[98]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[99], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[99]);
	$setuphold (posedge CPMFCMCLK, posedge FCMAPUSTOREDATA[9], 0:0:0, 0:0:0, notifier,,,CPMFCMCLK_delay,FCMAPUSTOREDATA_delay[9]);
	$setuphold (posedge CPMINTERCONNECTCLK, negedge CPMINTERCONNECTCLKNTO1, 0:0:0, 0:0:0, notifier,,,CPMINTERCONNECTCLK_delay,CPMINTERCONNECTCLKNTO1_delay);
	$setuphold (posedge CPMINTERCONNECTCLK, posedge CPMINTERCONNECTCLKNTO1, 0:0:0, 0:0:0, notifier,,,CPMINTERCONNECTCLK_delay,CPMINTERCONNECTCLKNTO1_delay);
	$setuphold (posedge CPMMCCLK, negedge MCMIADDRREADYTOACCEPT, 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIADDRREADYTOACCEPT_delay);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATAERR, 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATAERR_delay);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATAVALID, 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATAVALID_delay);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[0], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[0]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[100], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[100]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[101], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[101]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[102], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[102]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[103], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[103]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[104], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[104]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[105], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[105]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[106], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[106]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[107], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[107]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[108], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[108]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[109], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[109]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[10], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[10]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[110], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[110]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[111], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[111]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[112], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[112]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[113], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[113]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[114], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[114]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[115], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[115]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[116], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[116]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[117], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[117]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[118], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[118]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[119], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[119]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[11], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[11]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[120], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[120]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[121], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[121]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[122], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[122]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[123], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[123]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[124], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[124]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[125], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[125]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[126], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[126]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[127], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[127]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[12], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[12]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[13], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[13]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[14], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[14]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[15], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[15]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[16], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[16]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[17], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[17]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[18], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[18]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[19], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[19]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[1], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[1]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[20], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[20]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[21], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[21]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[22], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[22]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[23], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[23]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[24], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[24]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[25], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[25]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[26], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[26]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[27], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[27]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[28], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[28]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[29], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[29]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[2], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[2]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[30], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[30]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[31], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[31]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[32], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[32]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[33], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[33]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[34], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[34]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[35], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[35]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[36], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[36]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[37], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[37]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[38], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[38]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[39], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[39]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[3], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[3]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[40], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[40]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[41], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[41]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[42], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[42]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[43], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[43]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[44], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[44]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[45], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[45]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[46], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[46]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[47], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[47]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[48], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[48]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[49], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[49]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[4], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[4]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[50], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[50]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[51], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[51]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[52], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[52]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[53], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[53]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[54], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[54]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[55], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[55]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[56], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[56]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[57], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[57]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[58], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[58]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[59], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[59]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[5], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[5]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[60], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[60]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[61], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[61]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[62], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[62]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[63], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[63]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[64], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[64]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[65], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[65]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[66], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[66]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[67], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[67]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[68], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[68]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[69], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[69]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[6], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[6]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[70], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[70]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[71], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[71]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[72], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[72]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[73], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[73]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[74], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[74]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[75], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[75]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[76], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[76]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[77], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[77]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[78], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[78]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[79], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[79]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[7], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[7]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[80], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[80]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[81], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[81]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[82], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[82]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[83], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[83]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[84], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[84]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[85], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[85]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[86], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[86]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[87], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[87]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[88], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[88]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[89], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[89]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[8], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[8]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[90], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[90]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[91], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[91]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[92], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[92]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[93], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[93]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[94], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[94]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[95], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[95]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[96], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[96]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[97], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[97]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[98], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[98]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[99], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[99]);
	$setuphold (posedge CPMMCCLK, negedge MCMIREADDATA[9], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[9]);
	$setuphold (posedge CPMMCCLK, posedge MCMIADDRREADYTOACCEPT, 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIADDRREADYTOACCEPT_delay);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATAERR, 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATAERR_delay);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATAVALID, 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATAVALID_delay);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[0], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[0]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[100], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[100]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[101], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[101]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[102], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[102]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[103], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[103]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[104], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[104]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[105], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[105]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[106], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[106]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[107], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[107]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[108], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[108]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[109], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[109]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[10], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[10]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[110], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[110]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[111], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[111]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[112], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[112]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[113], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[113]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[114], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[114]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[115], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[115]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[116], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[116]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[117], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[117]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[118], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[118]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[119], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[119]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[11], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[11]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[120], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[120]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[121], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[121]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[122], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[122]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[123], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[123]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[124], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[124]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[125], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[125]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[126], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[126]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[127], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[127]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[12], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[12]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[13], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[13]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[14], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[14]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[15], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[15]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[16], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[16]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[17], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[17]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[18], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[18]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[19], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[19]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[1], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[1]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[20], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[20]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[21], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[21]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[22], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[22]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[23], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[23]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[24], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[24]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[25], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[25]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[26], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[26]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[27], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[27]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[28], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[28]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[29], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[29]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[2], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[2]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[30], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[30]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[31], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[31]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[32], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[32]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[33], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[33]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[34], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[34]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[35], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[35]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[36], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[36]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[37], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[37]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[38], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[38]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[39], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[39]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[3], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[3]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[40], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[40]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[41], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[41]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[42], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[42]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[43], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[43]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[44], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[44]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[45], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[45]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[46], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[46]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[47], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[47]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[48], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[48]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[49], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[49]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[4], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[4]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[50], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[50]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[51], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[51]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[52], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[52]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[53], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[53]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[54], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[54]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[55], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[55]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[56], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[56]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[57], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[57]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[58], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[58]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[59], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[59]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[5], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[5]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[60], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[60]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[61], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[61]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[62], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[62]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[63], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[63]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[64], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[64]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[65], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[65]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[66], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[66]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[67], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[67]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[68], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[68]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[69], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[69]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[6], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[6]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[70], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[70]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[71], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[71]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[72], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[72]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[73], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[73]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[74], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[74]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[75], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[75]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[76], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[76]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[77], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[77]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[78], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[78]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[79], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[79]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[7], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[7]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[80], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[80]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[81], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[81]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[82], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[82]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[83], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[83]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[84], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[84]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[85], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[85]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[86], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[86]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[87], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[87]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[88], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[88]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[89], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[89]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[8], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[8]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[90], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[90]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[91], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[91]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[92], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[92]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[93], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[93]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[94], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[94]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[95], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[95]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[96], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[96]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[97], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[97]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[98], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[98]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[99], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[99]);
	$setuphold (posedge CPMMCCLK, posedge MCMIREADDATA[9], 0:0:0, 0:0:0, notifier,,,CPMMCCLK_delay,MCMIREADDATA_delay[9]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMADDRACK, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMADDRACK_delay);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMMBUSY, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMMBUSY_delay);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMMIRQ, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMMIRQ_delay);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMMRDERR, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMMRDERR_delay);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMMWRERR, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMMWRERR_delay);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDBTERM, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDBTERM_delay);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDACK, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDACK_delay);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[0], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[0]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[100], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[100]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[101], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[101]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[102], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[102]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[103], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[103]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[104], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[104]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[105], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[105]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[106], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[106]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[107], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[107]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[108], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[108]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[109], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[109]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[10], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[10]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[110], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[110]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[111], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[111]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[112], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[112]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[113], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[113]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[114], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[114]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[115], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[115]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[116], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[116]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[117], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[117]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[118], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[118]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[119], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[119]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[11], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[11]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[120], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[120]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[121], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[121]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[122], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[122]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[123], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[123]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[124], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[124]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[125], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[125]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[126], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[126]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[127], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[127]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[12], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[12]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[13], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[13]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[14], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[14]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[15], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[15]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[16], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[16]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[17], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[17]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[18], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[18]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[19], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[19]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[1], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[1]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[20], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[20]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[21], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[21]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[22], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[22]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[23], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[23]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[24], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[24]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[25], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[25]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[26], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[26]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[27], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[27]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[28], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[28]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[29], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[29]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[2], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[2]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[30], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[30]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[31], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[31]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[32], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[32]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[33], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[33]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[34], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[34]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[35], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[35]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[36], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[36]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[37], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[37]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[38], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[38]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[39], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[39]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[3], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[3]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[40], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[40]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[41], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[41]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[42], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[42]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[43], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[43]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[44], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[44]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[45], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[45]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[46], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[46]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[47], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[47]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[48], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[48]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[49], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[49]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[4], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[4]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[50], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[50]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[51], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[51]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[52], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[52]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[53], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[53]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[54], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[54]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[55], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[55]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[56], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[56]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[57], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[57]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[58], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[58]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[59], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[59]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[5], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[5]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[60], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[60]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[61], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[61]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[62], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[62]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[63], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[63]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[64], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[64]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[65], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[65]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[66], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[66]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[67], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[67]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[68], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[68]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[69], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[69]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[6], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[6]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[70], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[70]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[71], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[71]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[72], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[72]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[73], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[73]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[74], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[74]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[75], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[75]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[76], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[76]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[77], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[77]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[78], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[78]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[79], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[79]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[7], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[7]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[80], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[80]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[81], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[81]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[82], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[82]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[83], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[83]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[84], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[84]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[85], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[85]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[86], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[86]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[87], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[87]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[88], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[88]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[89], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[89]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[8], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[8]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[90], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[90]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[91], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[91]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[92], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[92]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[93], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[93]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[94], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[94]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[95], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[95]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[96], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[96]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[97], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[97]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[98], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[98]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[99], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[99]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDDBUS[9], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[9]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDPENDPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDPENDPRI_delay[0]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDPENDPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDPENDPRI_delay[1]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDPENDREQ, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDPENDREQ_delay);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDWDADDR[0], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDWDADDR_delay[0]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDWDADDR[1], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDWDADDR_delay[1]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDWDADDR[2], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDWDADDR_delay[2]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMRDWDADDR[3], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDWDADDR_delay[3]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMREARBITRATE, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMREARBITRATE_delay);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMREQPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMREQPRI_delay[0]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMREQPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMREQPRI_delay[1]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMSSIZE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMSSIZE_delay[0]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMSSIZE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMSSIZE_delay[1]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMTIMEOUT, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMTIMEOUT_delay);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMWRBTERM, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMWRBTERM_delay);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMWRDACK, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMWRDACK_delay);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMWRPENDPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMWRPENDPRI_delay[0]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMWRPENDPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMWRPENDPRI_delay[1]);
	$setuphold (posedge CPMPPCMPLBCLK, negedge PLBPPCMWRPENDREQ, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMWRPENDREQ_delay);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMADDRACK, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMADDRACK_delay);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMMBUSY, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMMBUSY_delay);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMMIRQ, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMMIRQ_delay);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMMRDERR, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMMRDERR_delay);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMMWRERR, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMMWRERR_delay);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDBTERM, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDBTERM_delay);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDACK, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDACK_delay);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[0], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[0]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[100], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[100]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[101], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[101]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[102], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[102]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[103], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[103]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[104], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[104]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[105], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[105]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[106], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[106]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[107], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[107]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[108], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[108]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[109], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[109]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[10], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[10]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[110], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[110]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[111], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[111]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[112], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[112]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[113], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[113]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[114], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[114]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[115], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[115]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[116], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[116]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[117], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[117]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[118], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[118]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[119], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[119]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[11], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[11]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[120], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[120]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[121], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[121]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[122], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[122]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[123], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[123]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[124], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[124]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[125], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[125]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[126], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[126]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[127], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[127]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[12], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[12]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[13], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[13]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[14], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[14]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[15], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[15]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[16], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[16]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[17], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[17]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[18], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[18]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[19], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[19]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[1], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[1]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[20], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[20]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[21], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[21]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[22], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[22]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[23], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[23]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[24], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[24]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[25], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[25]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[26], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[26]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[27], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[27]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[28], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[28]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[29], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[29]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[2], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[2]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[30], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[30]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[31], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[31]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[32], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[32]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[33], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[33]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[34], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[34]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[35], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[35]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[36], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[36]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[37], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[37]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[38], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[38]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[39], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[39]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[3], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[3]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[40], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[40]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[41], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[41]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[42], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[42]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[43], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[43]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[44], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[44]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[45], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[45]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[46], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[46]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[47], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[47]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[48], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[48]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[49], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[49]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[4], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[4]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[50], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[50]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[51], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[51]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[52], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[52]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[53], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[53]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[54], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[54]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[55], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[55]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[56], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[56]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[57], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[57]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[58], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[58]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[59], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[59]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[5], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[5]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[60], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[60]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[61], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[61]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[62], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[62]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[63], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[63]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[64], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[64]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[65], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[65]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[66], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[66]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[67], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[67]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[68], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[68]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[69], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[69]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[6], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[6]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[70], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[70]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[71], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[71]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[72], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[72]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[73], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[73]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[74], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[74]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[75], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[75]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[76], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[76]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[77], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[77]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[78], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[78]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[79], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[79]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[7], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[7]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[80], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[80]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[81], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[81]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[82], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[82]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[83], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[83]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[84], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[84]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[85], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[85]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[86], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[86]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[87], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[87]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[88], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[88]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[89], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[89]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[8], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[8]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[90], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[90]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[91], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[91]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[92], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[92]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[93], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[93]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[94], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[94]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[95], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[95]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[96], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[96]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[97], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[97]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[98], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[98]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[99], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[99]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDDBUS[9], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDDBUS_delay[9]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDPENDPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDPENDPRI_delay[0]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDPENDPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDPENDPRI_delay[1]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDPENDREQ, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDPENDREQ_delay);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDWDADDR[0], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDWDADDR_delay[0]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDWDADDR[1], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDWDADDR_delay[1]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDWDADDR[2], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDWDADDR_delay[2]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMRDWDADDR[3], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMRDWDADDR_delay[3]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMREARBITRATE, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMREARBITRATE_delay);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMREQPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMREQPRI_delay[0]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMREQPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMREQPRI_delay[1]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMSSIZE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMSSIZE_delay[0]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMSSIZE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMSSIZE_delay[1]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMTIMEOUT, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMTIMEOUT_delay);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMWRBTERM, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMWRBTERM_delay);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMWRDACK, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMWRDACK_delay);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMWRPENDPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMWRPENDPRI_delay[0]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMWRPENDPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMWRPENDPRI_delay[1]);
	$setuphold (posedge CPMPPCMPLBCLK, posedge PLBPPCMWRPENDREQ, 0:0:0, 0:0:0, notifier,,,CPMPPCMPLBCLK_delay,PLBPPCMWRPENDREQ_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABORT, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABORT_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[10]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[11]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[12]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[13]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[14]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[15]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[16], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[16]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[17], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[17]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[18], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[18]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[19], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[19]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[20], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[20]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[21], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[21]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[22], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[22]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[23], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[23]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[24], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[24]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[25], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[25]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[26], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[26]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[27], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[27]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[28], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[28]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[29], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[29]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[2]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[30], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[30]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[31], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[31]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[3]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[4]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[5]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[6]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[7]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[8]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0ABUS[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[9]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[10]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[11]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[12]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[13]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[14]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[15]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[2]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[3]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[4]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[5]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[6]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[7]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[8]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BE[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[9]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0BUSLOCK, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BUSLOCK_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0LOCKERR, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0LOCKERR_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0MASTERID[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0MASTERID_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0MASTERID[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0MASTERID_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0MSIZE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0MSIZE_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0MSIZE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0MSIZE_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0PAVALID, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0PAVALID_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0RDBURST, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0RDBURST_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0RDPENDPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0RDPENDPRI_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0RDPENDPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0RDPENDPRI_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0RDPENDREQ, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0RDPENDREQ_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0RDPRIM, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0RDPRIM_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0REQPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0REQPRI_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0REQPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0REQPRI_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0RNW, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0RNW_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0SAVALID, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0SAVALID_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0SIZE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0SIZE_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0SIZE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0SIZE_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0SIZE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0SIZE_delay[2]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0SIZE[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0SIZE_delay[3]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[10]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[11]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[12]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[13]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[14]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[15]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[2]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[3]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[4]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[5]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[6]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[7]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[8]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TATTRIBUTE[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[9]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TYPE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TYPE_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TYPE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TYPE_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0TYPE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TYPE_delay[2]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0UABUS[28], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0UABUS_delay[28]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0UABUS[29], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0UABUS_delay[29]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0UABUS[30], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0UABUS_delay[30]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0UABUS[31], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0UABUS_delay[31]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRBURST, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRBURST_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[100], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[100]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[101], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[101]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[102], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[102]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[103], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[103]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[104], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[104]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[105], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[105]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[106], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[106]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[107], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[107]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[108], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[108]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[109], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[109]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[10]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[110], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[110]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[111], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[111]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[112], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[112]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[113], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[113]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[114], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[114]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[115], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[115]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[116], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[116]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[117], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[117]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[118], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[118]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[119], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[119]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[11]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[120], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[120]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[121], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[121]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[122], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[122]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[123], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[123]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[124], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[124]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[125], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[125]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[126], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[126]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[127], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[127]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[12]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[13]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[14]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[15]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[16], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[16]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[17], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[17]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[18], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[18]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[19], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[19]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[20], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[20]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[21], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[21]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[22], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[22]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[23], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[23]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[24], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[24]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[25], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[25]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[26], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[26]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[27], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[27]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[28], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[28]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[29], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[29]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[2]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[30], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[30]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[31], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[31]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[32], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[32]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[33], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[33]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[34], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[34]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[35], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[35]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[36], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[36]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[37], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[37]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[38], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[38]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[39], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[39]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[3]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[40], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[40]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[41], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[41]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[42], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[42]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[43], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[43]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[44], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[44]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[45], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[45]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[46], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[46]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[47], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[47]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[48], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[48]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[49], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[49]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[4]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[50], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[50]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[51], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[51]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[52], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[52]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[53], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[53]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[54], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[54]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[55], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[55]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[56], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[56]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[57], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[57]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[58], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[58]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[59], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[59]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[5]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[60], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[60]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[61], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[61]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[62], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[62]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[63], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[63]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[64], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[64]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[65], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[65]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[66], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[66]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[67], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[67]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[68], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[68]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[69], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[69]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[6]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[70], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[70]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[71], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[71]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[72], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[72]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[73], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[73]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[74], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[74]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[75], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[75]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[76], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[76]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[77], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[77]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[78], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[78]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[79], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[79]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[7]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[80], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[80]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[81], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[81]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[82], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[82]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[83], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[83]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[84], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[84]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[85], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[85]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[86], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[86]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[87], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[87]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[88], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[88]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[89], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[89]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[8]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[90], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[90]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[91], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[91]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[92], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[92]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[93], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[93]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[94], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[94]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[95], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[95]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[96], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[96]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[97], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[97]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[98], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[98]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[99], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[99]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRDBUS[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[9]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRPENDPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRPENDPRI_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRPENDPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRPENDPRI_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRPENDREQ, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRPENDREQ_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, negedge PLBPPCS0WRPRIM, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRPRIM_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABORT, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABORT_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[10]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[11]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[12]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[13]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[14]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[15]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[16], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[16]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[17], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[17]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[18], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[18]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[19], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[19]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[20], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[20]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[21], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[21]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[22], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[22]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[23], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[23]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[24], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[24]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[25], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[25]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[26], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[26]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[27], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[27]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[28], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[28]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[29], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[29]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[2]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[30], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[30]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[31], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[31]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[3]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[4]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[5]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[6]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[7]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[8]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0ABUS[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0ABUS_delay[9]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[10]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[11]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[12]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[13]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[14]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[15]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[2]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[3]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[4]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[5]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[6]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[7]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[8]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BE[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BE_delay[9]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0BUSLOCK, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0BUSLOCK_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0LOCKERR, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0LOCKERR_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0MASTERID[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0MASTERID_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0MASTERID[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0MASTERID_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0MSIZE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0MSIZE_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0MSIZE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0MSIZE_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0PAVALID, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0PAVALID_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0RDBURST, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0RDBURST_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0RDPENDPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0RDPENDPRI_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0RDPENDPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0RDPENDPRI_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0RDPENDREQ, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0RDPENDREQ_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0RDPRIM, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0RDPRIM_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0REQPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0REQPRI_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0REQPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0REQPRI_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0RNW, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0RNW_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0SAVALID, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0SAVALID_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0SIZE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0SIZE_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0SIZE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0SIZE_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0SIZE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0SIZE_delay[2]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0SIZE[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0SIZE_delay[3]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[10]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[11]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[12]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[13]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[14]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[15]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[2]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[3]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[4]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[5]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[6]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[7]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[8]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TATTRIBUTE[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TATTRIBUTE_delay[9]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TYPE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TYPE_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TYPE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TYPE_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0TYPE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0TYPE_delay[2]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0UABUS[28], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0UABUS_delay[28]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0UABUS[29], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0UABUS_delay[29]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0UABUS[30], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0UABUS_delay[30]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0UABUS[31], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0UABUS_delay[31]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRBURST, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRBURST_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[100], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[100]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[101], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[101]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[102], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[102]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[103], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[103]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[104], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[104]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[105], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[105]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[106], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[106]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[107], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[107]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[108], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[108]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[109], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[109]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[10]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[110], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[110]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[111], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[111]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[112], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[112]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[113], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[113]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[114], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[114]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[115], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[115]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[116], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[116]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[117], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[117]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[118], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[118]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[119], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[119]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[11]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[120], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[120]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[121], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[121]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[122], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[122]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[123], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[123]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[124], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[124]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[125], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[125]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[126], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[126]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[127], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[127]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[12]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[13]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[14]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[15]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[16], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[16]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[17], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[17]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[18], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[18]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[19], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[19]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[20], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[20]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[21], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[21]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[22], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[22]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[23], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[23]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[24], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[24]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[25], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[25]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[26], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[26]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[27], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[27]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[28], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[28]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[29], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[29]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[2]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[30], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[30]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[31], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[31]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[32], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[32]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[33], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[33]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[34], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[34]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[35], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[35]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[36], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[36]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[37], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[37]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[38], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[38]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[39], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[39]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[3]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[40], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[40]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[41], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[41]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[42], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[42]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[43], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[43]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[44], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[44]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[45], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[45]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[46], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[46]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[47], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[47]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[48], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[48]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[49], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[49]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[4]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[50], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[50]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[51], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[51]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[52], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[52]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[53], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[53]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[54], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[54]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[55], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[55]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[56], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[56]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[57], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[57]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[58], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[58]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[59], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[59]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[5]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[60], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[60]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[61], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[61]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[62], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[62]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[63], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[63]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[64], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[64]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[65], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[65]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[66], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[66]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[67], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[67]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[68], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[68]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[69], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[69]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[6]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[70], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[70]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[71], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[71]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[72], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[72]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[73], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[73]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[74], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[74]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[75], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[75]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[76], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[76]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[77], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[77]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[78], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[78]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[79], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[79]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[7]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[80], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[80]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[81], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[81]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[82], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[82]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[83], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[83]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[84], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[84]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[85], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[85]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[86], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[86]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[87], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[87]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[88], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[88]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[89], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[89]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[8]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[90], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[90]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[91], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[91]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[92], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[92]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[93], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[93]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[94], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[94]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[95], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[95]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[96], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[96]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[97], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[97]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[98], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[98]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[99], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[99]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRDBUS[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRDBUS_delay[9]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRPENDPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRPENDPRI_delay[0]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRPENDPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRPENDPRI_delay[1]);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRPENDREQ, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRPENDREQ_delay);
	$setuphold (posedge CPMPPCS0PLBCLK, posedge PLBPPCS0WRPRIM, 0:0:0, 0:0:0, notifier,,,CPMPPCS0PLBCLK_delay,PLBPPCS0WRPRIM_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABORT, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABORT_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[10]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[11]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[12]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[13]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[14]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[15]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[16], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[16]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[17], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[17]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[18], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[18]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[19], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[19]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[20], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[20]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[21], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[21]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[22], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[22]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[23], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[23]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[24], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[24]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[25], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[25]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[26], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[26]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[27], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[27]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[28], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[28]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[29], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[29]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[2]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[30], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[30]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[31], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[31]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[3]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[4]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[5]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[6]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[7]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[8]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1ABUS[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[9]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[10]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[11]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[12]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[13]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[14]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[15]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[2]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[3]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[4]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[5]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[6]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[7]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[8]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BE[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[9]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1BUSLOCK, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BUSLOCK_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1LOCKERR, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1LOCKERR_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1MASTERID[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1MASTERID_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1MASTERID[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1MASTERID_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1MSIZE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1MSIZE_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1MSIZE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1MSIZE_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1PAVALID, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1PAVALID_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1RDBURST, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1RDBURST_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1RDPENDPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1RDPENDPRI_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1RDPENDPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1RDPENDPRI_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1RDPENDREQ, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1RDPENDREQ_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1RDPRIM, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1RDPRIM_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1REQPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1REQPRI_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1REQPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1REQPRI_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1RNW, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1RNW_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1SAVALID, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1SAVALID_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1SIZE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1SIZE_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1SIZE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1SIZE_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1SIZE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1SIZE_delay[2]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1SIZE[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1SIZE_delay[3]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[10]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[11]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[12]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[13]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[14]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[15]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[2]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[3]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[4]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[5]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[6]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[7]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[8]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TATTRIBUTE[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[9]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TYPE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TYPE_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TYPE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TYPE_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1TYPE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TYPE_delay[2]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1UABUS[28], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1UABUS_delay[28]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1UABUS[29], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1UABUS_delay[29]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1UABUS[30], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1UABUS_delay[30]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1UABUS[31], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1UABUS_delay[31]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRBURST, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRBURST_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[100], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[100]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[101], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[101]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[102], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[102]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[103], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[103]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[104], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[104]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[105], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[105]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[106], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[106]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[107], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[107]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[108], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[108]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[109], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[109]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[10]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[110], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[110]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[111], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[111]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[112], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[112]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[113], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[113]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[114], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[114]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[115], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[115]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[116], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[116]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[117], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[117]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[118], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[118]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[119], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[119]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[11]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[120], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[120]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[121], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[121]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[122], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[122]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[123], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[123]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[124], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[124]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[125], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[125]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[126], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[126]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[127], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[127]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[12]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[13]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[14]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[15]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[16], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[16]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[17], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[17]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[18], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[18]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[19], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[19]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[20], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[20]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[21], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[21]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[22], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[22]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[23], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[23]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[24], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[24]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[25], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[25]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[26], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[26]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[27], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[27]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[28], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[28]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[29], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[29]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[2]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[30], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[30]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[31], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[31]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[32], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[32]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[33], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[33]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[34], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[34]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[35], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[35]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[36], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[36]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[37], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[37]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[38], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[38]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[39], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[39]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[3]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[40], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[40]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[41], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[41]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[42], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[42]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[43], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[43]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[44], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[44]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[45], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[45]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[46], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[46]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[47], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[47]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[48], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[48]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[49], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[49]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[4]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[50], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[50]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[51], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[51]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[52], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[52]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[53], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[53]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[54], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[54]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[55], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[55]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[56], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[56]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[57], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[57]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[58], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[58]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[59], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[59]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[5]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[60], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[60]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[61], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[61]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[62], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[62]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[63], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[63]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[64], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[64]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[65], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[65]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[66], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[66]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[67], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[67]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[68], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[68]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[69], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[69]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[6]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[70], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[70]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[71], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[71]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[72], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[72]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[73], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[73]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[74], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[74]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[75], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[75]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[76], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[76]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[77], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[77]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[78], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[78]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[79], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[79]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[7]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[80], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[80]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[81], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[81]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[82], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[82]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[83], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[83]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[84], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[84]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[85], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[85]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[86], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[86]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[87], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[87]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[88], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[88]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[89], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[89]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[8]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[90], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[90]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[91], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[91]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[92], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[92]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[93], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[93]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[94], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[94]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[95], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[95]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[96], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[96]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[97], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[97]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[98], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[98]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[99], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[99]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRDBUS[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[9]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRPENDPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRPENDPRI_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRPENDPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRPENDPRI_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRPENDREQ, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRPENDREQ_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, negedge PLBPPCS1WRPRIM, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRPRIM_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABORT, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABORT_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[10]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[11]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[12]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[13]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[14]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[15]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[16], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[16]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[17], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[17]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[18], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[18]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[19], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[19]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[20], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[20]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[21], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[21]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[22], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[22]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[23], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[23]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[24], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[24]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[25], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[25]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[26], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[26]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[27], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[27]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[28], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[28]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[29], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[29]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[2]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[30], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[30]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[31], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[31]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[3]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[4]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[5]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[6]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[7]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[8]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1ABUS[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1ABUS_delay[9]);  
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[10]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[11]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[12]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[13]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[14]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[15]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[2]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[3]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[4]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[5]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[6]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[7]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[8]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BE[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BE_delay[9]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1BUSLOCK, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1BUSLOCK_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1LOCKERR, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1LOCKERR_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1MASTERID[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1MASTERID_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1MASTERID[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1MASTERID_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1MSIZE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1MSIZE_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1MSIZE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1MSIZE_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1PAVALID, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1PAVALID_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1RDBURST, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1RDBURST_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1RDPENDPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1RDPENDPRI_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1RDPENDPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1RDPENDPRI_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1RDPENDREQ, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1RDPENDREQ_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1RDPRIM, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1RDPRIM_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1REQPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1REQPRI_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1REQPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1REQPRI_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1RNW, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1RNW_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1SAVALID, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1SAVALID_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1SIZE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1SIZE_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1SIZE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1SIZE_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1SIZE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1SIZE_delay[2]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1SIZE[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1SIZE_delay[3]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[10]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[11]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[12]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[13]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[14]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[15]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[2]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[3]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[4]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[5]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[6]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[7]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[8]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TATTRIBUTE[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TATTRIBUTE_delay[9]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TYPE[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TYPE_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TYPE[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TYPE_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1TYPE[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1TYPE_delay[2]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1UABUS[28], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1UABUS_delay[28]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1UABUS[29], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1UABUS_delay[29]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1UABUS[30], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1UABUS_delay[30]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1UABUS[31], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1UABUS_delay[31]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRBURST, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRBURST_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[100], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[100]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[101], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[101]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[102], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[102]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[103], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[103]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[104], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[104]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[105], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[105]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[106], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[106]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[107], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[107]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[108], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[108]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[109], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[109]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[10], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[10]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[110], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[110]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[111], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[111]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[112], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[112]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[113], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[113]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[114], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[114]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[115], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[115]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[116], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[116]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[117], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[117]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[118], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[118]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[119], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[119]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[11], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[11]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[120], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[120]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[121], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[121]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[122], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[122]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[123], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[123]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[124], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[124]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[125], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[125]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[126], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[126]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[127], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[127]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[12], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[12]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[13], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[13]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[14], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[14]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[15], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[15]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[16], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[16]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[17], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[17]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[18], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[18]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[19], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[19]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[20], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[20]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[21], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[21]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[22], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[22]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[23], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[23]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[24], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[24]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[25], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[25]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[26], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[26]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[27], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[27]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[28], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[28]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[29], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[29]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[2], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[2]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[30], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[30]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[31], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[31]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[32], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[32]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[33], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[33]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[34], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[34]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[35], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[35]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[36], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[36]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[37], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[37]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[38], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[38]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[39], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[39]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[3], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[3]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[40], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[40]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[41], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[41]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[42], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[42]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[43], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[43]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[44], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[44]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[45], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[45]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[46], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[46]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[47], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[47]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[48], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[48]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[49], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[49]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[4], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[4]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[50], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[50]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[51], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[51]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[52], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[52]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[53], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[53]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[54], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[54]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[55], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[55]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[56], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[56]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[57], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[57]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[58], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[58]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[59], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[59]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[5], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[5]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[60], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[60]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[61], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[61]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[62], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[62]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[63], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[63]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[64], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[64]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[65], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[65]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[66], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[66]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[67], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[67]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[68], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[68]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[69], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[69]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[6], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[6]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[70], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[70]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[71], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[71]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[72], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[72]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[73], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[73]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[74], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[74]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[75], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[75]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[76], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[76]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[77], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[77]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[78], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[78]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[79], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[79]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[7], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[7]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[80], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[80]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[81], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[81]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[82], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[82]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[83], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[83]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[84], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[84]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[85], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[85]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[86], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[86]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[87], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[87]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[88], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[88]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[89], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[89]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[8], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[8]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[90], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[90]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[91], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[91]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[92], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[92]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[93], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[93]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[94], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[94]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[95], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[95]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[96], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[96]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[97], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[97]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[98], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[98]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[99], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[99]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRDBUS[9], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRDBUS_delay[9]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRPENDPRI[0], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRPENDPRI_delay[0]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRPENDPRI[1], 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRPENDPRI_delay[1]);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRPENDREQ, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRPENDREQ_delay);
	$setuphold (posedge CPMPPCS1PLBCLK, posedge PLBPPCS1WRPRIM, 0:0:0, 0:0:0, notifier,,,CPMPPCS1PLBCLK_delay,PLBPPCS1WRPRIM_delay);
	$setuphold (posedge JTGC440TCK, negedge CPMC440CORECLOCKINACTIVE, 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,CPMC440CORECLOCKINACTIVE_delay);
	$setuphold (posedge JTGC440TCK, negedge DBGC440SYSTEMSTATUS[0], 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,DBGC440SYSTEMSTATUS_delay[0]);
	$setuphold (posedge JTGC440TCK, negedge DBGC440SYSTEMSTATUS[1], 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,DBGC440SYSTEMSTATUS_delay[1]);
	$setuphold (posedge JTGC440TCK, negedge DBGC440SYSTEMSTATUS[2], 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,DBGC440SYSTEMSTATUS_delay[2]);
	$setuphold (posedge JTGC440TCK, negedge DBGC440SYSTEMSTATUS[3], 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,DBGC440SYSTEMSTATUS_delay[3]);
	$setuphold (posedge JTGC440TCK, negedge DBGC440SYSTEMSTATUS[4], 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,DBGC440SYSTEMSTATUS_delay[4]);
	$setuphold (posedge JTGC440TCK, negedge JTGC440TDI, 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,JTGC440TDI_delay);
	$setuphold (posedge JTGC440TCK, negedge JTGC440TMS, 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,JTGC440TMS_delay);
	$setuphold (posedge JTGC440TCK, posedge CPMC440CORECLOCKINACTIVE, 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,CPMC440CORECLOCKINACTIVE_delay);
	$setuphold (posedge JTGC440TCK, posedge DBGC440SYSTEMSTATUS[0], 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,DBGC440SYSTEMSTATUS_delay[0]);
	$setuphold (posedge JTGC440TCK, posedge DBGC440SYSTEMSTATUS[1], 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,DBGC440SYSTEMSTATUS_delay[1]);
	$setuphold (posedge JTGC440TCK, posedge DBGC440SYSTEMSTATUS[2], 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,DBGC440SYSTEMSTATUS_delay[2]);
	$setuphold (posedge JTGC440TCK, posedge DBGC440SYSTEMSTATUS[3], 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,DBGC440SYSTEMSTATUS_delay[3]);
	$setuphold (posedge JTGC440TCK, posedge DBGC440SYSTEMSTATUS[4], 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,DBGC440SYSTEMSTATUS_delay[4]);
	$setuphold (posedge JTGC440TCK, posedge JTGC440TDI, 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,JTGC440TDI_delay);
	$setuphold (posedge JTGC440TCK, posedge JTGC440TMS, 0:0:0, 0:0:0, notifier,,,JTGC440TCK_delay,JTGC440TMS_delay);
	(CPMC440CLK => C440CPMCORESLEEPREQ) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440CPMDECIRPTREQ) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440CPMFITIRPTREQ) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440CPMMSRCE) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440CPMMSREE) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440CPMTIMERRESETREQ) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440CPMWDIRPTREQ) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440DBGSYSTEMCONTROL[0]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440DBGSYSTEMCONTROL[1]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440DBGSYSTEMCONTROL[2]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440DBGSYSTEMCONTROL[3]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440DBGSYSTEMCONTROL[4]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440DBGSYSTEMCONTROL[5]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440DBGSYSTEMCONTROL[6]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440DBGSYSTEMCONTROL[7]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440MACHINECHECK) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCBRANCHSTATUS[0]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCBRANCHSTATUS[1]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCBRANCHSTATUS[2]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCCYCLE) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCEXECUTIONSTATUS[0]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCEXECUTIONSTATUS[1]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCEXECUTIONSTATUS[2]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCEXECUTIONSTATUS[3]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCEXECUTIONSTATUS[4]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRACESTATUS[0]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRACESTATUS[1]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRACESTATUS[2]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRACESTATUS[3]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRACESTATUS[4]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRACESTATUS[5]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRACESTATUS[6]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTOUT) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE[0]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE[10]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE[11]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE[12]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE[13]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE[1]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE[2]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE[3]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE[4]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE[5]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE[6]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE[7]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE[8]) = (100:100:100, 100:100:100);
	(CPMC440CLK => C440TRCTRIGGEREVENTTYPE[9]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRABUS[0]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRABUS[1]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRABUS[2]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRABUS[3]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRABUS[4]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRABUS[5]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRABUS[6]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRABUS[7]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRABUS[8]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRABUS[9]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[0]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[10]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[11]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[12]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[13]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[14]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[15]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[16]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[17]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[18]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[19]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[1]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[20]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[21]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[22]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[23]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[24]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[25]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[26]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[27]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[28]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[29]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[2]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[30]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[31]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[3]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[4]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[5]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[6]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[7]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[8]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRDBUSOUT[9]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRREAD) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRUABUS[20]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRUABUS[21]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDMDCRWRITE) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRACK) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[0]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[10]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[11]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[12]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[13]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[14]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[15]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[16]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[17]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[18]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[19]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[1]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[20]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[21]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[22]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[23]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[24]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[25]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[26]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[27]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[28]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[29]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[2]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[30]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[31]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[3]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[4]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[5]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[6]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[7]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[8]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRDBUSIN[9]) = (100:100:100, 100:100:100);
	(CPMDCRCLK => PPCDSDCRTIMEOUTWAIT) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLRSTENGINEACK) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLRXDSTRDYN) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[0]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[10]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[11]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[12]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[13]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[14]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[15]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[16]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[17]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[18]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[19]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[1]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[20]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[21]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[22]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[23]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[24]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[25]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[26]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[27]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[28]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[29]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[2]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[30]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[31]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[3]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[4]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[5]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[6]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[7]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[8]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXD[9]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXEOFN) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXEOPN) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXREM[0]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXREM[1]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXREM[2]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXREM[3]) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXSOFN) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXSOPN) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0LLTXSRCRDYN) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0RXIRQ) = (100:100:100, 100:100:100);
	(CPMDMA0LLCLK => DMA0TXIRQ) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLRSTENGINEACK) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLRXDSTRDYN) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[0]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[10]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[11]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[12]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[13]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[14]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[15]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[16]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[17]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[18]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[19]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[1]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[20]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[21]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[22]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[23]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[24]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[25]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[26]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[27]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[28]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[29]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[2]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[30]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[31]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[3]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[4]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[5]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[6]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[7]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[8]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXD[9]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXEOFN) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXEOPN) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXREM[0]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXREM[1]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXREM[2]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXREM[3]) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXSOFN) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXSOPN) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1LLTXSRCRDYN) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1RXIRQ) = (100:100:100, 100:100:100);
	(CPMDMA1LLCLK => DMA1TXIRQ) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLRSTENGINEACK) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLRXDSTRDYN) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[0]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[10]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[11]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[12]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[13]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[14]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[15]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[16]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[17]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[18]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[19]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[1]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[20]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[21]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[22]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[23]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[24]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[25]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[26]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[27]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[28]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[29]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[2]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[30]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[31]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[3]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[4]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[5]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[6]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[7]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[8]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXD[9]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXEOFN) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXEOPN) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXREM[0]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXREM[1]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXREM[2]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXREM[3]) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXSOFN) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXSOPN) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2LLTXSRCRDYN) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2RXIRQ) = (100:100:100, 100:100:100);
	(CPMDMA2LLCLK => DMA2TXIRQ) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLRSTENGINEACK) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLRXDSTRDYN) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[0]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[10]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[11]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[12]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[13]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[14]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[15]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[16]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[17]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[18]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[19]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[1]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[20]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[21]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[22]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[23]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[24]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[25]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[26]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[27]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[28]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[29]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[2]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[30]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[31]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[3]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[4]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[5]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[6]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[7]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[8]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXD[9]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXEOFN) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXEOPN) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXREM[0]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXREM[1]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXREM[2]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXREM[3]) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXSOFN) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXSOPN) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3LLTXSRCRDYN) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3RXIRQ) = (100:100:100, 100:100:100);
	(CPMDMA3LLCLK => DMA3TXIRQ) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMDECFPUOP) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMDECLDSTXFERSIZE[0]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMDECLDSTXFERSIZE[1]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMDECLDSTXFERSIZE[2]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMDECLOAD) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMDECNONAUTON) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMDECSTORE) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMDECUDIVALID) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMDECUDI[0]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMDECUDI[1]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMDECUDI[2]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMDECUDI[3]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMENDIAN) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMFLUSH) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[0]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[10]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[11]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[12]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[13]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[14]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[15]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[16]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[17]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[18]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[19]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[1]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[20]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[21]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[22]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[23]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[24]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[25]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[26]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[27]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[28]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[29]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[2]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[30]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[31]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[3]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[4]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[5]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[6]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[7]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[8]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRUCTION[9]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMINSTRVALID) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADBYTEADDR[0]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADBYTEADDR[1]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADBYTEADDR[2]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADBYTEADDR[3]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[0]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[100]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[101]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[102]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[103]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[104]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[105]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[106]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[107]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[108]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[109]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[10]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[110]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[111]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[112]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[113]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[114]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[115]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[116]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[117]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[118]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[119]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[11]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[120]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[121]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[122]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[123]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[124]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[125]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[126]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[127]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[12]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[13]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[14]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[15]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[16]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[17]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[18]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[19]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[1]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[20]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[21]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[22]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[23]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[24]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[25]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[26]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[27]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[28]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[29]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[2]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[30]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[31]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[32]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[33]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[34]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[35]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[36]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[37]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[38]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[39]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[3]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[40]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[41]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[42]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[43]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[44]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[45]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[46]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[47]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[48]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[49]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[4]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[50]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[51]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[52]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[53]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[54]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[55]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[56]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[57]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[58]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[59]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[5]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[60]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[61]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[62]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[63]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[64]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[65]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[66]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[67]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[68]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[69]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[6]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[70]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[71]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[72]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[73]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[74]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[75]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[76]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[77]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[78]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[79]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[7]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[80]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[81]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[82]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[83]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[84]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[85]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[86]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[87]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[88]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[89]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[8]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[90]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[91]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[92]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[93]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[94]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[95]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[96]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[97]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[98]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[99]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDATA[9]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMLOADDVALID) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMMSRFE0) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMMSRFE1) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMNEXTINSTRREADY) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMOPERANDVALID) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[0]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[10]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[11]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[12]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[13]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[14]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[15]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[16]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[17]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[18]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[19]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[1]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[20]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[21]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[22]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[23]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[24]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[25]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[26]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[27]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[28]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[29]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[2]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[30]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[31]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[3]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[4]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[5]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[6]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[7]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[8]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRADATA[9]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[0]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[10]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[11]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[12]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[13]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[14]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[15]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[16]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[17]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[18]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[19]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[1]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[20]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[21]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[22]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[23]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[24]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[25]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[26]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[27]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[28]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[29]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[2]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[30]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[31]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[3]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[4]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[5]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[6]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[7]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[8]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMRBDATA[9]) = (100:100:100, 100:100:100);
	(CPMFCMCLK => APUFCMWRITEBACKOK) = (100:100:100, 100:100:100);
	(CPMINTERCONNECTCLK => C440RSTCHIPRESETREQ) = (100:100:100, 100:100:100);
	(CPMINTERCONNECTCLK => C440RSTCORERESETREQ) = (100:100:100, 100:100:100);
	(CPMINTERCONNECTCLK => C440RSTSYSTEMRESETREQ) = (100:100:100, 100:100:100);
	(CPMINTERCONNECTCLK => PPCCPMINTERCONNECTBUSY) = (100:100:100, 100:100:100);
	(CPMINTERCONNECTCLK => PPCEICINTERCONNECTIRQ) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESSVALID) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[0]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[10]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[11]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[12]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[13]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[14]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[15]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[16]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[17]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[18]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[19]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[1]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[20]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[21]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[22]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[23]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[24]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[25]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[26]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[27]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[28]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[29]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[2]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[30]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[31]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[32]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[33]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[34]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[35]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[3]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[4]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[5]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[6]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[7]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[8]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCADDRESS[9]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBANKCONFLICT) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[0]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[10]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[11]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[12]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[13]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[14]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[15]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[1]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[2]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[3]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[4]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[5]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[6]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[7]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[8]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCBYTEENABLE[9]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCREADNOTWRITE) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCROWCONFLICT) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATAVALID) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[0]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[100]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[101]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[102]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[103]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[104]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[105]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[106]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[107]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[108]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[109]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[10]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[110]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[111]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[112]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[113]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[114]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[115]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[116]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[117]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[118]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[119]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[11]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[120]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[121]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[122]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[123]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[124]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[125]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[126]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[127]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[12]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[13]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[14]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[15]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[16]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[17]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[18]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[19]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[1]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[20]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[21]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[22]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[23]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[24]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[25]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[26]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[27]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[28]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[29]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[2]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[30]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[31]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[32]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[33]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[34]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[35]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[36]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[37]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[38]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[39]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[3]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[40]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[41]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[42]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[43]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[44]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[45]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[46]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[47]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[48]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[49]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[4]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[50]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[51]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[52]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[53]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[54]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[55]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[56]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[57]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[58]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[59]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[5]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[60]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[61]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[62]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[63]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[64]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[65]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[66]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[67]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[68]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[69]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[6]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[70]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[71]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[72]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[73]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[74]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[75]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[76]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[77]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[78]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[79]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[7]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[80]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[81]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[82]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[83]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[84]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[85]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[86]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[87]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[88]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[89]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[8]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[90]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[91]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[92]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[93]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[94]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[95]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[96]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[97]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[98]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[99]) = (100:100:100, 100:100:100);
	(CPMMCCLK => MIMCWRITEDATA[9]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABORT) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[0]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[10]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[11]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[12]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[13]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[14]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[15]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[16]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[17]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[18]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[19]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[1]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[20]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[21]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[22]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[23]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[24]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[25]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[26]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[27]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[28]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[29]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[2]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[30]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[31]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[3]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[4]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[5]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[6]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[7]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[8]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBABUS[9]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[0]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[10]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[11]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[12]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[13]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[14]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[15]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[1]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[2]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[3]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[4]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[5]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[6]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[7]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[8]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBE[9]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBBUSLOCK) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBLOCKERR) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBPRIORITY[0]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBPRIORITY[1]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBRDBURST) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBREQUEST) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBRNW) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBSIZE[0]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBSIZE[1]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBSIZE[2]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBSIZE[3]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[0]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[10]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[11]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[12]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[13]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[14]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[15]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[1]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[2]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[3]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[4]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[5]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[6]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[7]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[8]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTATTRIBUTE[9]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTYPE[0]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTYPE[1]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBTYPE[2]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBUABUS[28]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBUABUS[29]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBUABUS[30]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBUABUS[31]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRBURST) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[0]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[100]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[101]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[102]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[103]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[104]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[105]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[106]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[107]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[108]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[109]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[10]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[110]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[111]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[112]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[113]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[114]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[115]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[116]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[117]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[118]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[119]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[11]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[120]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[121]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[122]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[123]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[124]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[125]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[126]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[127]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[12]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[13]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[14]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[15]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[16]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[17]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[18]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[19]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[1]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[20]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[21]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[22]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[23]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[24]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[25]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[26]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[27]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[28]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[29]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[2]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[30]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[31]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[32]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[33]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[34]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[35]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[36]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[37]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[38]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[39]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[3]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[40]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[41]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[42]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[43]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[44]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[45]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[46]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[47]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[48]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[49]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[4]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[50]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[51]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[52]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[53]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[54]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[55]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[56]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[57]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[58]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[59]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[5]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[60]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[61]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[62]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[63]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[64]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[65]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[66]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[67]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[68]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[69]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[6]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[70]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[71]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[72]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[73]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[74]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[75]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[76]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[77]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[78]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[79]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[7]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[80]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[81]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[82]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[83]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[84]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[85]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[86]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[87]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[88]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[89]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[8]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[90]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[91]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[92]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[93]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[94]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[95]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[96]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[97]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[98]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[99]) = (100:100:100, 100:100:100);
	(CPMPPCMPLBCLK => PPCMPLBWRDBUS[9]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBADDRACK) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMBUSY[0]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMBUSY[1]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMBUSY[2]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMBUSY[3]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMIRQ[0]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMIRQ[1]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMIRQ[2]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMIRQ[3]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMRDERR[0]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMRDERR[1]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMRDERR[2]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMRDERR[3]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMWRERR[0]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMWRERR[1]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMWRERR[2]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBMWRERR[3]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDBTERM) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDCOMP) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDACK) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[0]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[100]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[101]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[102]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[103]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[104]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[105]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[106]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[107]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[108]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[109]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[10]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[110]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[111]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[112]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[113]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[114]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[115]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[116]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[117]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[118]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[119]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[11]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[120]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[121]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[122]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[123]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[124]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[125]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[126]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[127]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[12]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[13]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[14]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[15]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[16]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[17]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[18]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[19]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[1]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[20]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[21]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[22]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[23]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[24]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[25]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[26]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[27]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[28]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[29]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[2]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[30]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[31]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[32]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[33]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[34]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[35]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[36]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[37]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[38]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[39]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[3]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[40]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[41]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[42]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[43]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[44]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[45]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[46]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[47]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[48]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[49]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[4]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[50]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[51]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[52]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[53]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[54]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[55]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[56]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[57]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[58]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[59]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[5]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[60]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[61]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[62]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[63]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[64]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[65]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[66]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[67]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[68]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[69]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[6]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[70]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[71]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[72]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[73]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[74]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[75]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[76]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[77]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[78]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[79]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[7]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[80]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[81]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[82]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[83]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[84]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[85]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[86]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[87]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[88]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[89]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[8]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[90]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[91]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[92]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[93]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[94]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[95]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[96]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[97]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[98]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[99]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDDBUS[9]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDWDADDR[0]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDWDADDR[1]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDWDADDR[2]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBRDWDADDR[3]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBREARBITRATE) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBSSIZE[0]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBSSIZE[1]) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBWAIT) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBWRBTERM) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBWRCOMP) = (100:100:100, 100:100:100);
	(CPMPPCS0PLBCLK => PPCS0PLBWRDACK) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBADDRACK) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMBUSY[0]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMBUSY[1]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMBUSY[2]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMBUSY[3]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMIRQ[0]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMIRQ[1]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMIRQ[2]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMIRQ[3]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMRDERR[0]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMRDERR[1]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMRDERR[2]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMRDERR[3]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMWRERR[0]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMWRERR[1]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMWRERR[2]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBMWRERR[3]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDBTERM) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDCOMP) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDACK) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[0]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[100]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[101]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[102]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[103]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[104]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[105]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[106]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[107]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[108]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[109]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[10]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[110]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[111]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[112]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[113]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[114]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[115]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[116]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[117]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[118]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[119]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[11]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[120]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[121]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[122]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[123]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[124]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[125]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[126]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[127]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[12]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[13]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[14]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[15]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[16]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[17]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[18]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[19]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[1]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[20]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[21]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[22]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[23]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[24]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[25]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[26]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[27]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[28]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[29]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[2]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[30]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[31]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[32]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[33]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[34]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[35]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[36]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[37]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[38]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[39]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[3]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[40]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[41]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[42]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[43]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[44]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[45]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[46]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[47]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[48]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[49]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[4]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[50]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[51]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[52]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[53]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[54]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[55]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[56]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[57]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[58]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[59]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[5]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[60]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[61]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[62]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[63]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[64]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[65]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[66]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[67]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[68]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[69]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[6]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[70]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[71]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[72]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[73]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[74]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[75]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[76]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[77]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[78]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[79]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[7]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[80]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[81]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[82]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[83]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[84]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[85]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[86]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[87]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[88]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[89]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[8]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[90]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[91]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[92]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[93]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[94]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[95]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[96]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[97]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[98]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[99]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDDBUS[9]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDWDADDR[0]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDWDADDR[1]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDWDADDR[2]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBRDWDADDR[3]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBREARBITRATE) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBSSIZE[0]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBSSIZE[1]) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBWAIT) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBWRBTERM) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBWRCOMP) = (100:100:100, 100:100:100);
	(CPMPPCS1PLBCLK => PPCS1PLBWRDACK) = (100:100:100, 100:100:100);
	(JTGC440TCK => C440JTGTDO) = (100:100:100, 100:100:100);
	(JTGC440TCK => C440JTGTDOEN) = (100:100:100, 100:100:100);

	specparam PATHPULSE$ = 0;
endspecify
endmodule
