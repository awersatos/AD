--------------------------------------------------------------------
--       Actel A500K VITAL Library
--       NAME: a500k.vhd
--       DATE: May 17, 2006
---------------------------------------------------------------------/



library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.VITAL_Timing.all;

package COMPONENTS is

constant DefaultTimingChecksOn : Boolean := True;
constant DefaultXGenerationOn : Boolean := False;
constant DefaultXon : Boolean := False;
constant DefaultMsgOn : Boolean := True;



------ Component AND2 ------
 component AND2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND2FT ------
 component AND2FT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND3 ------
 component AND3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND3FFT ------
 component AND3FFT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AND3FTT ------
 component AND3FTT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO21 ------
 component AO21
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO21FTF ------
 component AO21FTF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO21FTT ------
 component AO21FTT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AO21TTF ------
 component AO21TTF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI21 ------
 component AOI21
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI21FTF ------
 component AOI21FTF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI21FTT ------
 component AOI21FTT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component AOI21TTF ------
 component AOI21TTF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BFR ------
 component BFR
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component BUBBLE ------
 component BUBBLE
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component DMUX ------
 component DMUX
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component GL25 ------
 component GL25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GL25LP ------
 component GL25LP
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GL25LPU ------
 component GL25LPU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GL25U ------
 component GL25U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GL33 ------
 component GL33
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GL33U ------
 component GL33U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLINT ------
 component GLINT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GND ------
 component GND
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True		);
    port(
		Y		: out    STD_ULOGIC);
 end component;


------ Component IB25 ------
 component IB25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IB25LP ------
 component IB25LP
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IB25LPU ------
 component IB25LPU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IB25U ------
 component IB25U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IB33 ------
 component IB33
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IB33U ------
 component IB33U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component INV ------
 component INV
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component LD ------
 component LD
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component LDB ------
 component LDB
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component LDBI ------
 component LDBI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component LDC ------
 component LDC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component LDCI ------
 component LDCI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component LDI ------
 component LDI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component LDL ------
 component LDL
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component LDLB ------
 component LDLB
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component LDLBI ------
 component LDLBI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component LDLC ------
 component LDLC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component LDLCI ------
 component LDLCI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component LDLI ------
 component LDLI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component LDLS ------
 component LDLS
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component LDLSI ------
 component LDLSI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component LDS ------
 component LDS
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component LDSI ------
 component LDSI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component MUX2H ------
 component MUX2H
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component MUX2L ------
 component MUX2L
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND2 ------
 component NAND2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND2FT ------
 component NAND2FT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND3 ------
 component NAND3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND3FFT ------
 component NAND3FFT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NAND3FTT ------
 component NAND3FTT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR2 ------
 component NOR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR2FT ------
 component NOR2FT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR3 ------
 component NOR3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR3FFT ------
 component NOR3FFT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NOR3FTT ------
 component NOR3FTT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component NUBBLE ------
 component NUBBLE
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA21 ------
 component OA21
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA21FTF ------
 component OA21FTF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA21FTT ------
 component OA21FTT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OA21TTF ------
 component OA21TTF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OAI21 ------
 component OAI21
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OAI21FTF ------
 component OAI21FTF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OAI21FTT ------
 component OAI21FTT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OAI21TTF ------
 component OAI21TTF
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		C		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OB25HH ------
 component OB25HH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB25HL ------
 component OB25HL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB25HN ------
 component OB25HN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB25LH ------
 component OB25LH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB25LL ------
 component OB25LL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB25LN ------
 component OB25LN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB25LPHH ------
 component OB25LPHH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB25LPHL ------
 component OB25LPHL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB25LPHN ------
 component OB25LPHN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB25LPLH ------
 component OB25LPLH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB25LPLL ------
 component OB25LPLL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB25LPLN ------
 component OB25LPLN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB33LH ------
 component OB33LH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB33LL ------
 component OB33LL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB33LN ------
 component OB33LN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB33PH ------
 component OB33PH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB33PL ------
 component OB33PL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OB33PN ------
 component OB33PN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OR2 ------
 component OR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR2FT ------
 component OR2FT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR3 ------
 component OR3
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR3FFT ------
 component OR3FFT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OR3FTT ------
 component OR3FTT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component PWR ------
 component PWR
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True		);
    port(
		Y		: out    STD_ULOGIC);
 end component;


------ Component XNOR2 ------
 component XNOR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XNOR2FT ------
 component XNOR2FT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XOR2 ------
 component XOR2
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component XOR2FT ------
 component XOR2FT
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component DFF ------
 component DFF
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFFB ------
 component DFFB
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFFBI ------
 component DFFBI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component DFFC ------
 component DFFC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFFCI ------
 component DFFCI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component DFFI ------
 component DFFI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component DFFL ------
 component DFFL
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFFLB ------
 component DFFLB
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFFLBI ------
 component DFFLBI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component DFFLC ------
 component DFFLC
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFFLCI ------
 component DFFLCI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component DFFLI ------
 component DFFLI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component DFFLS ------
 component DFFLS
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFFLSI ------
 component DFFLSI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component DFFS ------
 component DFFS
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 end component;


------ Component DFFSI ------
 component DFFSI
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 end component;


------ Component GLIB25 ------
 component GLIB25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLIB25LP ------
 component GLIB25LP
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLIB25LPU ------
 component GLIB25LPU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLIB25U ------
 component GLIB25U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLIB33 ------
 component GLIB33
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLIB33U ------
 component GLIB33U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLMIB25 ------
 component GLMIB25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLMIB33 ------
 component GLMIB33
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLMIB25LP ------
 component GLMIB25LP
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLMIB25U ------
 component GLMIB25U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLMIB33U ------
 component GLMIB33U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLMIB25LPU ------
 component GLMIB25LPU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLMIBL25 ------
 component GLMIBL25
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLMIBL33 ------
 component GLMIBL33
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLMIBL25LP ------
 component GLMIBL25LP
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLMIBL25LPU ------
 component GLMIBL25LPU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLMIBL33U ------
 component GLMIBL33U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component GLMIBL25U ------
 component GLMIBL25U
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 end component;


------ Component IOB25HH ------
 component IOB25HH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
       		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25HL ------
 component IOB25HL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25HN ------
 component IOB25HN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LH ------
 component IOB25LH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LL ------
 component IOB25LL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
                tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LN ------
 component IOB25LN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25HHU ------
 component IOB25HHU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25HLU ------
 component IOB25HLU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25HNU ------
 component IOB25HNU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LHU ------
 component IOB25LHU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LLU ------
 component IOB25LLU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LNU ------
 component IOB25LNU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LPHH ------
 component IOB25LPHH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LPHL ------
 component IOB25LPHL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LPHN ------
 component IOB25LPHN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LPLH ------
 component IOB25LPLH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LPLL ------
 component IOB25LPLL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LPLN ------
 component IOB25LPLN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LPHHU ------
 component IOB25LPHHU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LPHLU ------
 component IOB25LPHLU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LPHNU ------
 component IOB25LPHNU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LPLHU ------
 component IOB25LPLHU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LPLLU ------
 component IOB25LPLLU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB25LPLNU ------
 component IOB25LPLNU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB33LH ------
 component IOB33LH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB33LL ------
 component IOB33LL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB33LN ------
 component IOB33LN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB33PH ------
 component IOB33PH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB33PL ------
 component IOB33PL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB33PN ------
 component IOB33PN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB33LHU ------
 component IOB33LHU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB33LLU ------
 component IOB33LLU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB33LNU ------
 component IOB33LNU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB33PHU ------
 component IOB33PHU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB33PLU ------
 component IOB33PLU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOB33PNU ------
 component IOB33PNU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25HH ------
 component IOBL25HH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25HL ------
 component IOBL25HL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25HN ------
 component IOBL25HN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LH ------
 component IOBL25LH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LL ------
 component IOBL25LL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LN ------
 component IOBL25LN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25HHU ------
 component IOBL25HHU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25HLU ------
 component IOBL25HLU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25HNU ------
 component IOBL25HNU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LHU ------
 component IOBL25LHU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LLU ------
 component IOBL25LLU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LNU ------
 component IOBL25LNU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LPHH ------
 component IOBL25LPHH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LPHL ------
 component IOBL25LPHL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LPHN ------
 component IOBL25LPHN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LPLH ------
 component IOBL25LPLH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LPLL ------
 component IOBL25LPLL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LPLN ------
 component IOBL25LPLN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LPHHU ------
 component IOBL25LPHHU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LPHLU ------
 component IOBL25LPHLU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LPHNU ------
 component IOBL25LPHNU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LPLHU ------
 component IOBL25LPLHU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LPLLU ------
 component IOBL25LPLLU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL25LPLNU ------
 component IOBL25LPLNU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL33LH ------
 component IOBL33LH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL33LL ------
 component IOBL33LL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL33LN ------
 component IOBL33LN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL33PH ------
 component IOBL33PH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL33PL ------
 component IOBL33PL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL33PN ------
 component IOBL33PN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL33LHU ------
 component IOBL33LHU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL33LLU ------
 component IOBL33LLU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL33LNU ------
 component IOBL33LNU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL33PHU ------
 component IOBL33PHU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL33PLU ------
 component IOBL33PLU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component IOBL33PNU ------
 component IOBL33PNU
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 end component;


------ Component OTB25HH ------
 component OTB25HH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB25HL ------
 component OTB25HL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB25HN ------
 component OTB25HN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB25LH ------
 component OTB25LH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB25LL ------
 component OTB25LL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB25LN ------
 component OTB25LN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB25LPLH ------
 component OTB25LPLH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB25LPLL ------
 component OTB25LPLL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB25LPLN ------
 component OTB25LPLN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB25LPHH ------
 component OTB25LPHH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB25LPHL ------
 component OTB25LPHL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB25LPHN ------
 component OTB25LPHN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB33LH ------
 component OTB33LH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB33LL ------
 component OTB33LL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB33LN ------
 component OTB33LN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB33PH ------
 component OTB33PH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB33PL ------
 component OTB33PL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTB33PN ------
 component OTB33PN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL25HH ------
 component OTBL25HH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL25HL ------
 component OTBL25HL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL25HN ------
 component OTBL25HN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL25LH ------
 component OTBL25LH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL25LL ------
 component OTBL25LL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL25LN ------
 component OTBL25LN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL25LPLH ------
 component OTBL25LPLH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL25LPLL ------
 component OTBL25LPLL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL25LPLN ------
 component OTBL25LPLN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL25LPHH ------
 component OTBL25LPHH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL25LPHL ------
 component OTBL25LPHL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL25LPHN ------
 component OTBL25LPHN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL33LH ------
 component OTBL33LH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL33LL ------
 component OTBL33LL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL33LN ------
 component OTBL33LN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL33PH ------
 component OTBL33PH
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL33PL ------
 component OTBL33PL
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;


------ Component OTBL33PN ------
 component OTBL33PN
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 end component;

component RAM256x9AA
   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI0_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI1_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI2_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI3_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI4_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI5_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI6_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI7_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI8_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns,0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpw_RDB_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_RDB_negedge	        : VitalDelayType := 0.000 ns;
 	tperiod_RDB	        : VitalDelayType := 0.000 ns;
 	tpw_RBLKB_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RBLKB_negedge	: VitalDelayType := 0.000 ns;
 	tperiod_RBLKB	        : VitalDelayType := 0.000 ns;
 	tpw_RADDR0_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR0_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                           : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                         : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                         : VitalDelayType := 0.000 ns;
 	tperiod_WRB                             : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_RDB_WRB_negedge_negedge          : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_WRB_posedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RBLKB_WRB_posedge_posedge         : VitalDelayType := 0.000 ns;
 	thold_RDB_WBLKB_posedge_posedge         : VitalDelayType := 0.000 ns;
 	thold_RBLKB_WBLKB_posedge_posedge       : VitalDelayType := 0.000 ns;
 	thold_RADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';
   WPE    :  OUT STD_LOGIC := 'X';
   RPE    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');
end component;

component RAM256x9AAP
   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpw_RDB_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_RDB_negedge	        : VitalDelayType := 0.000 ns;
 	tperiod_RDB	        : VitalDelayType := 0.000 ns;
 	tpw_RBLKB_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RBLKB_negedge	: VitalDelayType := 0.000 ns;
 	tperiod_RBLKB	        : VitalDelayType := 0.000 ns;
 	tpw_RADDR0_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR0_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                           : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                         : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                         : VitalDelayType := 0.000 ns;
 	tperiod_WRB                             : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_RDB_WRB_negedge_negedge          : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_WRB_posedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RBLKB_WRB_posedge_posedge         : VitalDelayType := 0.000 ns;
 	thold_RDB_WBLKB_posedge_posedge         : VitalDelayType := 0.000 ns;
 	thold_RBLKB_WBLKB_posedge_posedge       : VitalDelayType := 0.000 ns;
 	thold_RADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');
end component;

component RAM256x9AST
   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI0_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI1_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI2_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI3_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI4_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI5_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI6_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI7_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI8_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                           : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                         : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                         : VitalDelayType := 0.000 ns;
 	tperiod_WRB                             : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WRB_RCLKS_negedge_posedge        : VitalDelayType := 0.000 ns;
 	thold_WRB_RCLKS_negedge_posedge         : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RCLKS_negedge_posedge      : VitalDelayType := 0.000 ns;
	thold_WBLKB_RCLKS_negedge_posedge       : VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';
   WPE    :  OUT STD_LOGIC := 'X';
   RPE    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');
end component;

component RAM256x9ASTP
   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                           : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                         : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                         : VitalDelayType := 0.000 ns;
 	tperiod_WRB                             : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WRB_RCLKS_negedge_posedge        : VitalDelayType := 0.000 ns;
 	thold_WRB_RCLKS_negedge_posedge         : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RCLKS_negedge_posedge      : VitalDelayType := 0.000 ns;
	thold_WBLKB_RCLKS_negedge_posedge       : VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');
end component;

component RAM256x9ASR
   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI0_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI1_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI2_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI3_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI4_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI5_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI6_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI7_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI8_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                           : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                         : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                         : VitalDelayType := 0.000 ns;
 	tperiod_WRB                             : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WRB_RCLKS_negedge_posedge        : VitalDelayType := 0.000 ns;
 	thold_WRB_RCLKS_negedge_posedge         : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RCLKS_negedge_posedge      : VitalDelayType := 0.000 ns;
	thold_WBLKB_RCLKS_negedge_posedge       : VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';
   WPE    :  OUT STD_LOGIC := 'X';
   RPE    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');
end component;

component RAM256x9ASRP
   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                           : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                         : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                         : VitalDelayType := 0.000 ns;
 	tperiod_WRB                             : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WRB_RCLKS_negedge_posedge        : VitalDelayType := 0.000 ns;
 	thold_WRB_RCLKS_negedge_posedge         : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RCLKS_negedge_posedge      : VitalDelayType := 0.000 ns;
	thold_WBLKB_RCLKS_negedge_posedge       : VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');
end component;

component RAM256x9SA
   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_WCLKS_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns,0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpw_RDB_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_RDB_negedge	        : VitalDelayType := 0.000 ns;
 	tperiod_RDB	        : VitalDelayType := 0.000 ns;
 	tpw_RBLKB_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RBLKB_negedge	: VitalDelayType := 0.000 ns;
 	tperiod_RBLKB	        : VitalDelayType := 0.000 ns;
 	tpw_RADDR0_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR0_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tpw_WCLKS_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                           : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_RDB_WCLKS_negedge_posedge       : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_WCLKS_negedge_posedge       : VitalDelayType := 0.000 ns;
 	tsetup_RADDR0_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR0_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR1_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR2_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR3_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR4_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR5_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR6_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR7_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	thold_RDB_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RBLKB_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR0_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR1_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR2_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR3_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR4_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR5_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR6_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR7_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';
   WPE    :  OUT STD_LOGIC := 'X';
   RPE    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   WCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');
end component;

component RAM256x9SAP
   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpw_RDB_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_RDB_negedge	        : VitalDelayType := 0.000 ns;
 	tperiod_RDB	        : VitalDelayType := 0.000 ns;
 	tpw_RBLKB_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RBLKB_negedge	: VitalDelayType := 0.000 ns;
 	tperiod_RBLKB	        : VitalDelayType := 0.000 ns;
 	tpw_RADDR0_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR0_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tpw_WCLKS_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                           : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_RDB_WCLKS_negedge_posedge       : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_WCLKS_negedge_posedge       : VitalDelayType := 0.000 ns;
 	tsetup_RADDR0_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR0_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR1_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR2_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR3_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR4_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR5_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR6_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR7_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	thold_RDB_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RBLKB_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR0_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR1_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR2_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR3_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR4_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR5_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR6_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR7_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   WCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');
end component;

component RAM256x9SST
   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_WCLKS_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tpw_WCLKS_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                           : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 7.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';
   WPE    :  OUT STD_LOGIC := 'X';
   RPE    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   WCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');
end component;

component RAM256x9SSTP
   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tpw_WCLKS_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                           : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 7.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   WCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');
end component;

component RAM256x9SSR
   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_WCLKS_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tpw_WCLKS_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                           : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 7.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';
   WPE    :  OUT STD_LOGIC := 'X';
   RPE    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   WCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');
end component;

component RAM256x9SSRP
   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tpw_WCLKS_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                           : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 7.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   WCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');
end component;


component FIFO256x9AA
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI0_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI1_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI2_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI3_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI4_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI5_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI6_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI7_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI8_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tpw_RDB_posedge         : VitalDelayType        := 0.000 ns;
 	tpw_RDB_negedge         : VitalDelayType        := 0.000 ns;
 	tperiod_RDB             : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_posedge       : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_negedge       : VitalDelayType        := 0.000 ns;
 	tperiod_RBLKB           : VitalDelayType        := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;

  	-- WB falling edge hold to RESETB   
 	thold_WRB_RESET_posedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_RESET_posedge_posedge             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_RESET_posedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RESET_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_WRB_RESET_negedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WBLKB_RESET_negedge_posedge             : VitalDelayType := 0.000 ns;
	tsetup_WRB_RESET_negedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_RESET_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                               : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                               : VitalDelayType := 0.000 ns;
 	tperiod_WRB                                   : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        WPE    :  OUT STD_LOGIC := 'X';
        RPE    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');

end component;

component FIFO256x9AAP
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tpw_RDB_posedge         : VitalDelayType        := 0.000 ns;
 	tpw_RDB_negedge         : VitalDelayType        := 0.000 ns;
 	tperiod_RDB             : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_posedge       : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_negedge       : VitalDelayType        := 0.000 ns;
 	tperiod_RBLKB           : VitalDelayType        := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;

  	-- WB falling edge hold to RESETB   
 	thold_WRB_RESET_posedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_RESET_posedge_posedge             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_RESET_posedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RESET_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_WRB_RESET_negedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WBLKB_RESET_negedge_posedge             : VitalDelayType := 0.000 ns;
	tsetup_WRB_RESET_negedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_RESET_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                               : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                               : VitalDelayType := 0.000 ns;
 	tperiod_WRB                                   : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');

end component;

component FIFO256x9AST
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI0_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI1_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI2_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI3_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI4_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI5_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI6_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI7_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI8_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;

  	-- WB falling edge hold to RESETB   
 	thold_WRB_RESET_posedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_RESET_posedge_posedge             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_RESET_posedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RESET_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_WRB_RESET_negedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WBLKB_RESET_negedge_posedge             : VitalDelayType := 0.000 ns;
	tsetup_WRB_RESET_negedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_RESET_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                               : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                               : VitalDelayType := 0.000 ns;
 	tperiod_WRB                                   : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        WPE    :  OUT STD_LOGIC := 'X';
        RPE    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');

end component;

component FIFO256x9ASTP
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;

  	-- WB falling edge hold to RESETB   
 	thold_WRB_RESET_posedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_RESET_posedge_posedge             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_RESET_posedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RESET_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_WRB_RESET_negedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WBLKB_RESET_negedge_posedge             : VitalDelayType := 0.000 ns;
	tsetup_WRB_RESET_negedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_RESET_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                               : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                               : VitalDelayType := 0.000 ns;
 	tperiod_WRB                                   : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');

end component;

component FIFO256x9ASR
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI0_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI1_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI2_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI3_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI4_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI5_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI6_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI7_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI8_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;

  	-- WB falling edge hold to RESETB   
 	thold_WRB_RESET_posedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_RESET_posedge_posedge             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_RESET_posedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RESET_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_WRB_RESET_negedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WBLKB_RESET_negedge_posedge             : VitalDelayType := 0.000 ns;
	tsetup_WRB_RESET_negedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_RESET_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                               : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                               : VitalDelayType := 0.000 ns;
 	tperiod_WRB                                   : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        WPE    :  OUT STD_LOGIC := 'X';
        RPE    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');

end component;

component FIFO256x9ASRP
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;

  	-- WB falling edge hold to RESETB   
 	thold_WRB_RESET_posedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_RESET_posedge_posedge             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_RESET_posedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RESET_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_WRB_RESET_negedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WBLKB_RESET_negedge_posedge             : VitalDelayType := 0.000 ns;
	tsetup_WRB_RESET_negedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_RESET_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                               : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                               : VitalDelayType := 0.000 ns;
 	tperiod_WRB                                   : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');

end component;

component FIFO256x9SA
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_PARODD_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tpw_RDB_posedge         : VitalDelayType        := 0.000 ns;
 	tpw_RDB_negedge         : VitalDelayType        := 0.000 ns;
 	tperiod_RDB             : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_posedge       : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_negedge       : VitalDelayType        := 0.000 ns;
 	tperiod_RBLKB           : VitalDelayType        := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_WCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_WCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;

        -- WCLK falling edge setup to RESET rising edge 
 	trecovery_RESET_WCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_WCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- WCLK rising  edge hold to RESET rising edge 
	thold_RESET_WCLKS_posedge_posedge             : VitalDelayType := 0.00 ns;
	thold_RESET_WCLKS_posedge_negedge             : VitalDelayType := 0.00 ns;
	tpw_WCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        WPE    :  OUT STD_LOGIC := 'X';
        RPE    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        WCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');

end component;

component FIFO256x9SAP
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tpw_RDB_posedge         : VitalDelayType        := 0.000 ns;
 	tpw_RDB_negedge         : VitalDelayType        := 0.000 ns;
 	tperiod_RDB             : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_posedge       : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_negedge       : VitalDelayType        := 0.000 ns;
 	tperiod_RBLKB           : VitalDelayType        := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_WCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_WCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;

        -- WCLK falling edge setup to RESET rising edge 
 	trecovery_RESET_WCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_WCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- WCLK rising  edge hold to RESET rising edge 
	thold_RESET_WCLKS_posedge_posedge             : VitalDelayType := 0.00 ns;
	thold_RESET_WCLKS_posedge_negedge             : VitalDelayType := 0.00 ns;
	tpw_WCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        WCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');

end component;

component FIFO256x9SST
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_PARODD_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_WCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_WCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;

        -- WCLK falling edge setup to RESET rising edge 
 	trecovery_RESET_WCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_WCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- WCLK rising  edge hold to RESET rising edge 
	thold_RESET_WCLKS_posedge_posedge             : VitalDelayType := 0.00 ns;
	thold_RESET_WCLKS_posedge_negedge             : VitalDelayType := 0.00 ns;
	tpw_WCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        WPE    :  OUT STD_LOGIC := 'X';
        RPE    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        WCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');

end component;

component FIFO256x9SSTP
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_WCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_WCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;

        -- WCLK falling edge setup to RESET rising edge 
 	trecovery_RESET_WCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_WCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- WCLK rising  edge hold to RESET rising edge 
	thold_RESET_WCLKS_posedge_posedge             : VitalDelayType := 0.00 ns;
	thold_RESET_WCLKS_posedge_negedge             : VitalDelayType := 0.00 ns;
	tpw_WCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        WCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');

end component;

component FIFO256x9SSR
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_PARODD_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_WCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_WCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;

        -- WCLK falling edge setup to RESET rising edge 
 	trecovery_RESET_WCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_WCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- WCLK rising  edge hold to RESET rising edge 
	thold_RESET_WCLKS_posedge_posedge             : VitalDelayType := 0.00 ns;
	thold_RESET_WCLKS_posedge_negedge             : VitalDelayType := 0.00 ns;
	tpw_WCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        WPE    :  OUT STD_LOGIC := 'X';
        RPE    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        WCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');

end component;

component FIFO256x9SSRP
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_WCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_WCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;

        -- WCLK falling edge setup to RESET rising edge 
 	trecovery_RESET_WCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_WCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- WCLK rising  edge hold to RESET rising edge 
	thold_RESET_WCLKS_posedge_posedge             : VitalDelayType := 0.00 ns;
	thold_RESET_WCLKS_posedge_negedge             : VitalDelayType := 0.00 ns;
	tpw_WCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        WCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');

end component;

component UJTAG
      generic(
      tipd_UTDO      : VitalDelayType01 := (  0.0 ns,0.0 ns );
      tipd_TMS       : VitalDelayType01 := (  0.0 ns,0.0 ns );
      tipd_TDI       : VitalDelayType01 := (  0.0 ns,0.0 ns );
      tipd_TCK       : VitalDelayType01 := (  0.0 ns,0.0 ns );
      tipd_TRSTB     : VitalDelayType01 := (  0.0 ns,0.0 ns );

      TimingChecksOn : Boolean := True;
      InstancePath   : String  := "*";
      Xon            : Boolean := False;
      MsgOn          : Boolean := True);

    port(
      UTDO           :  in    STD_ULOGIC;
      TMS            :  in    STD_ULOGIC;
      TDI            :  in    STD_ULOGIC;
      TCK            :  in    STD_ULOGIC;
      TRSTB          :  in    STD_ULOGIC;
      UIREG0         :  out   STD_ULOGIC;
      UIREG1         :  out   STD_ULOGIC;
      UIREG2         :  out   STD_ULOGIC;
      UIREG3         :  out   STD_ULOGIC;
      UIREG4         :  out   STD_ULOGIC;
      UIREG5         :  out   STD_ULOGIC;
      UIREG6         :  out   STD_ULOGIC;
      UIREG7         :  out   STD_ULOGIC;
      UTDI           :  out   STD_ULOGIC;
      URSTB          :  out   STD_ULOGIC;
      UDRCK          :  out   STD_ULOGIC;
      UDRSH          :  out   STD_ULOGIC;
      UDRUPD         :  out   STD_ULOGIC;
      TDO            :  out   STD_ULOGIC);
end component;

end COMPONENTS;

--------------------- END OF COMPONENTS PACKAGE SECTION  ----------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;

use IEEE.VITAL_Timing.all;
use IEEE.VITAL_Primitives.all;

package VTABLES is

   CONSTANT L : VitalTableSymbolType := '0';
   CONSTANT H : VitalTableSymbolType := '1';
   CONSTANT x : VitalTableSymbolType := '-';
   CONSTANT S : VitalTableSymbolType := 'S';
   CONSTANT R : VitalTableSymbolType := '/';
   CONSTANT U : VitalTableSymbolType := 'X';
   CONSTANT V : VitalTableSymbolType := 'B'; -- valid clock signal (non-rising)

-- CLR_ipd, CLK_delayed, Q_zd, D, E_delayed, PRE_ipd, CLK_ipd
CONSTANT DFEG_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  x,  x,  x,  L ),
( H,  L,  H,  H,  x,  x,  H,  x,  H ),
( H,  L,  H,  x,  H,  x,  H,  x,  H ),
( H,  L,  x,  H,  L,  x,  H,  x,  H ),
( H,  H,  x,  x,  x,  H,  x,  x,  S ),
( H,  x,  x,  x,  x,  L,  x,  x,  H ),
( H,  x,  x,  x,  x,  H,  L,  x,  S ),
( x,  L,  L,  L,  x,  H,  H,  x,  L ),
( x,  L,  L,  x,  H,  H,  H,  x,  L ),
( x,  L,  x,  L,  L,  H,  H,  x,  L ),
( U,  x,  L,  x,  x,  H,  x,  x,  L ),
( H,  x,  H,  x,  x,  U,  x,  x,  H )); 

-- CLR_ipd, CLK_delayed, T_delayed, Q_zd, CLK_ipd
CONSTANT tflipflop_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  x,  L ),
( H,  L,  L,  H,  H,  x,  H ),
( H,  L,  H,  L,  H,  x,  H ),
( H,  H,  x,  x,  x,  x,  S ),
( H,  x,  x,  x,  L,  x,  S ),
( x,  L,  L,  L,  H,  x,  L ),
( x,  L,  H,  H,  H,  x,  L ));

-- CLR_ipd, CLK_delayed, PRE_delayed,K_delayed,J_delayed, Q_zd, CLK_ipd
CONSTANT jkflipflop_Q_tab : VitalStateTableType := (
( L,  x,  H,  x,  x,  x,  x,  x,  U ),
( L,  x,  L,  x,  x,  x,  x,  x,  L ),
( H,  L,  x,  L,  H,  x,  H,  x,  H ),
( H,  L,  x,  L,  x,  H,  H,  x,  H ),
( H,  L,  x,  x,  H,  L,  H,  x,  H ),
( H,  H,  L,  x,  x,  x,  x,  x,  S ),
( H,  x,  L,  x,  x,  x,  L,  x,  S ),
( H,  x,  H,  x,  x,  x,  x,  x,  H ),
( x,  L,  L,  H,  L,  x,  H,  x,  L ),
( x,  L,  L,  H,  x,  H,  H,  x,  L ),
( x,  L,  L,  x,  L,  L,  H,  x,  L ),
( U,  x,  L,  x,  x,  L,  x,  x,  L ),
( H,  x,  U,  x,  x,  H,  x,  x,  H ));

CONSTANT JKF2A_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  x,  x,  L ),
( H,  L,  L,  H,  x,  H,  x,  H ),
( H,  L,  L,  x,  H,  H,  x,  H ),
( H,  L,  x,  H,  L,  H,  x,  H ),
( H,  H,  x,  x,  x,  x,  x,  S ),
( H,  x,  x,  x,  x,  L,  x,  S ),
( x,  L,  H,  L,  x,  H,  x,  L ),
( x,  L,  H,  x,  H,  H,  x,  L ),
( x,  L,  x,  L,  L,  H,  x,  L ),
( U,  x,  x,  x,  L,  x,  x,  L ));

CONSTANT JKF3A_Q_tab : VitalStateTableType := (
( L,  H,  L,  x,  H,  H,  x,  L ),
( L,  H,  x,  H,  H,  H,  x,  L ),
( L,  L,  H,  x,  x,  H,  x,  H ),
( L,  L,  x,  H,  x,  H,  x,  H ),
( L,  x,  L,  L,  H,  H,  x,  L ),
( L,  x,  H,  L,  x,  H,  x,  H ),
( H,  x,  x,  x,  H,  x,  x,  S ),
( x,  x,  x,  x,  L,  x,  x,  H ),
( x,  x,  x,  x,  H,  L,  x,  S ),
( x,  x,  x,  H,  U,  x,  x,  H ));

CONSTANT dlatch_DLE3B_Q_tab : VitalStateTableType := (
( x,  x,  x,  H,  x,  H ),   --active high preset

( H,  x,  x,  L,  x,  S ),   --latch
( x,  H,  x,  L,  x,  S ),   --latch

( L,  L,  H,  L,  x,  H ),   --transparent
( L,  L,  L,  L,  x,  L ),   --transparent

( U,  x,  H,  L,  H,  H ),   --o/p mux pessimism
( x,  U,  H,  L,  H,  H ),   --o/p mux pessimism
( U,  x,  L,  L,  L,  L ),   --o/p mux pessimism
( x,  U,  L,  L,  L,  L ),   --o/p mux pessimism

( L,  L,  H,  U,  x,  H ),   --PRE==X
( H,  x,  x,  U,  H,  H ),   --PRE==X
( x,  H,  x,  U,  H,  H ),   --PRE==X
( L,  U,  H,  U,  H,  H ),   --PRE==X
( U,  L,  H,  U,  H,  H ),   --PRE==X
( U,  U,  H,  U,  H,  H ));  --PRE==X
--G, E, D, P, Qn, Qn+1

CONSTANT dlatch_DLE2B_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  L ),   --active low clear

( H,  H,  x,  x,  x,  S ),   --latch
( H,  x,  H,  x,  x,  S ),   --latch

( H,  L,  L,  H,  x,  H ),   --transparent
( H,  L,  L,  L,  x,  L ),   --transparent

( H,  x,  x,  L,  L,  L ),   --o/p mux pessimism
( H,  x,  x,  H,  H,  H ),   --o/p mux pessimism

( U,  x,  x,  L,  L,  L ),   --CLR==X, o/p mux pessimism
( U,  H,  x,  x,  L,  L ),   --CLR==X, o/p mux pessimism, latch
( U,  x,  H,  x,  L,  L ),   --CLR==X, o/p mux pessimism, latch
( U,  L,  L,  L,  x,  L ));  --CLR==X, i/p mux pessimism
--C, G, E, D, Qn, Qn+1


CONSTANT dlatch_DL2C_Q_tab : VitalStateTableType := (
( L,  x,  x,  x,  x,  L ),   --active low clear
( H,  x,  x,  H,  x,  H ),   --active high preset

( H,  H,  x,  L,  x,  S ),   --latch
( H,  L,  L,  L,  x,  L ),   --transparent

( U,  L,  L,  L,  x,  L ),   --CLR==U
( U,  H,  x,  L,  L,  L ),   --CLR==U
( x,  U,  L,  L,  L,  L ),   --CLR,G==U

( H,  U,  H,  x,  H,  H ),   --PRE==U/x,G==U
( H,  L,  H,  x,  x,  H ),   --PRE==U/x
( H,  H,  x,  U,  H,  H ));  --PRE==U
--CLR, G, D, PRE, Qn, Qn+1

end VTABLES;



--------------------- END OF VITABLE TABLE SECTION  ----------------



 ---- CELL AND2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND2 :  entity is True;
 end AND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of AND2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( A_ipd  AND  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND2_VITAL of AND2 is 
    for VITAL_ACT
    end for;
 end CFG_AND2_VITAL;



 ---- CELL AND2FT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND2FT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND2FT :  entity is True;
 end AND2FT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of AND2FT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT A_ipd)  AND  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND2FT_VITAL of AND2FT is 
    for VITAL_ACT
    end for;
 end CFG_AND2FT_VITAL;



 ---- CELL AND3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND3 :  entity is True;
 end AND3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of AND3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND3_VITAL of AND3 is 
    for VITAL_ACT
    end for;
 end CFG_AND3_VITAL;



 ---- CELL AND3FFT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND3FFT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND3FFT :  entity is True;
 end AND3FFT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of AND3FFT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND3FFT_VITAL of AND3FFT is 
    for VITAL_ACT
    end for;
 end CFG_AND3FFT_VITAL;



 ---- CELL AND3FTT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AND3FTT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AND3FTT :  entity is True;
 end AND3FTT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of AND3FTT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  B_ipd ) AND  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AND3FTT_VITAL of AND3FTT is 
    for VITAL_ACT
    end for;
 end CFG_AND3FTT_VITAL;



 ---- CELL AO21 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO21 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO21 :  entity is True;
 end AO21;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of AO21 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO21_VITAL of AO21 is 
    for VITAL_ACT
    end for;
 end CFG_AO21_VITAL;



 ---- CELL AO21FTF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO21FTF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO21FTF :  entity is True;
 end AO21FTF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of AO21FTF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  B_ipd ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO21FTF_VITAL of AO21FTF is 
    for VITAL_ACT
    end for;
 end CFG_AO21FTF_VITAL;



 ---- CELL AO21FTT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO21FTT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO21FTT :  entity is True;
 end AO21FTT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of AO21FTT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO21FTT_VITAL of AO21FTT is 
    for VITAL_ACT
    end for;
 end CFG_AO21FTT_VITAL;



 ---- CELL AO21TTF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AO21TTF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AO21TTF :  entity is True;
 end AO21TTF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of AO21TTF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AO21TTF_VITAL of AO21TTF is 
    for VITAL_ACT
    end for;
 end CFG_AO21TTF_VITAL;



 ---- CELL AOI21 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI21 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI21 :  entity is True;
 end AOI21;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of AOI21 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, C_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT C_ipd) ) OR ( (NOT B_ipd)  AND  (NOT C_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (C_ipd'last_event,tpd_C_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI21_VITAL of AOI21 is 
    for VITAL_ACT
    end for;
 end CFG_AOI21_VITAL;



 ---- CELL AOI21FTF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI21FTF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI21FTF :  entity is True;
 end AOI21FTF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of AOI21FTF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, C_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  C_ipd ) OR ( (NOT B_ipd)  AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (C_ipd'last_event,tpd_C_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI21FTF_VITAL of AOI21FTF is 
    for VITAL_ACT
    end for;
 end CFG_AOI21FTF_VITAL;



 ---- CELL AOI21FTT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI21FTT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI21FTT :  entity is True;
 end AOI21FTT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of AOI21FTT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, C_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  (NOT C_ipd) ) OR ( (NOT B_ipd)  AND  (NOT C_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (C_ipd'last_event,tpd_C_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI21FTT_VITAL of AOI21FTT is 
    for VITAL_ACT
    end for;
 end CFG_AOI21FTT_VITAL;



 ---- CELL AOI21TTF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity AOI21TTF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of AOI21TTF :  entity is True;
 end AOI21TTF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of AOI21TTF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, C_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  C_ipd ) OR ( (NOT B_ipd)  AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (C_ipd'last_event,tpd_C_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_AOI21TTF_VITAL of AOI21TTF is 
    for VITAL_ACT
    end for;
 end CFG_AOI21TTF_VITAL;



 ---- CELL BFR ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BFR is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BFR :  entity is True;
 end BFR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of BFR is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BFR_VITAL of BFR is 
    for VITAL_ACT
    end for;
 end CFG_BFR_VITAL;



 ---- CELL BUBBLE ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity BUBBLE is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of BUBBLE :  entity is True;
 end BUBBLE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of BUBBLE is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  (NOT A_ipd) ;


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_BUBBLE_VITAL of BUBBLE is 
    for VITAL_ACT
    end for;
 end CFG_BUBBLE_VITAL;



 ---- CELL DMUX ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DMUX is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of DMUX :  entity is True;
 end DMUX;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DMUX is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (S_ipd'last_event,tpd_S_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_DMUX_VITAL of DMUX is 
    for VITAL_ACT
    end for;
 end CFG_DMUX_VITAL;



 ---- CELL GL25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GL25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GL25 :  entity is True;
 end GL25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GL25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS GL_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        GL_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GL25_VITAL of GL25 is 
    for VITAL_ACT
    end for;
 end CFG_GL25_VITAL;



 ---- CELL GL25LP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GL25LP is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GL25LP :  entity is True;
 end GL25LP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GL25LP is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS GL_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        GL_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GL25LP_VITAL of GL25LP is 
    for VITAL_ACT
    end for;
 end CFG_GL25LP_VITAL;



 ---- CELL GL25LPU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GL25LPU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GL25LPU :  entity is True;
 end GL25LPU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GL25LPU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS GL_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        GL_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GL25LPU_VITAL of GL25LPU is 
    for VITAL_ACT
    end for;
 end CFG_GL25LPU_VITAL;



 ---- CELL GL25U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GL25U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GL25U :  entity is True;
 end GL25U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GL25U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS GL_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        GL_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GL25U_VITAL of GL25U is 
    for VITAL_ACT
    end for;
 end CFG_GL25U_VITAL;



 ---- CELL GL33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GL33 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GL33 :  entity is True;
 end GL33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GL33 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS GL_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        GL_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GL33_VITAL of GL33 is 
    for VITAL_ACT
    end for;
 end CFG_GL33_VITAL;



 ---- CELL GL33U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GL33U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GL33U :  entity is True;
 end GL33U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GL33U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS GL_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        GL_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GL33U_VITAL of GL33U is 
    for VITAL_ACT
    end for;
 end CFG_GL33U_VITAL;



 ---- CELL GLINT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLINT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLINT :  entity is True;
 end GLINT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLINT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS GL_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        GL_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLINT_VITAL of GLINT is 
    for VITAL_ACT
    end for;
 end CFG_GLINT_VITAL;



 ---- CELL GND ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GND is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True		);
    port(
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GND :  entity is True;
 end GND;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GND is
	attribute VITAL_LEVEL0 of VITAL_ACT : architecture is True;


begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	--- Empty
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
        Y<= '0';


end VITAL_ACT;

 configuration CFG_GND_VITAL of GND is 
    for VITAL_ACT
    end for;
 end CFG_GND_VITAL;



 ---- CELL IB25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IB25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IB25 :  entity is True;
 end IB25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IB25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IB25_VITAL of IB25 is 
    for VITAL_ACT
    end for;
 end CFG_IB25_VITAL;



 ---- CELL IB25LP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IB25LP is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IB25LP :  entity is True;
 end IB25LP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IB25LP is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IB25LP_VITAL of IB25LP is 
    for VITAL_ACT
    end for;
 end CFG_IB25LP_VITAL;



 ---- CELL IB25LPU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IB25LPU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IB25LPU :  entity is True;
 end IB25LPU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IB25LPU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IB25LPU_VITAL of IB25LPU is 
    for VITAL_ACT
    end for;
 end CFG_IB25LPU_VITAL;



 ---- CELL IB25U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IB25U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IB25U :  entity is True;
 end IB25U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IB25U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IB25U_VITAL of IB25U is 
    for VITAL_ACT
    end for;
 end CFG_IB25U_VITAL;



 ---- CELL IB33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IB33 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IB33 :  entity is True;
 end IB33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IB33 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IB33_VITAL of IB33 is 
    for VITAL_ACT
    end for;
 end CFG_IB33_VITAL;



 ---- CELL IB33U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IB33U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IB33U :  entity is True;
 end IB33U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IB33U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IB33U_VITAL of IB33U is 
    for VITAL_ACT
    end for;
 end CFG_IB33U_VITAL;



 ---- CELL INV ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity INV is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of INV :  entity is True;
 end INV;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of INV is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  (NOT A_ipd) ;


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_INV_VITAL of INV is 
    for VITAL_ACT
    end for;
 end CFG_INV_VITAL;



 ---- CELL LD ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LD is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LD :  entity is True;
 end LD;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LD is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_negedge,
	 TimingData		=> Tmkr_D_EN_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_negedge,
	 SetupLow		=> tsetup_D_EN_negedge_negedge,
	 HoldHigh		=> thold_D_EN_posedge_negedge,
	 HoldLow		=> thold_D_EN_negedge_negedge,
	 CheckEnabled		=>  True, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/LD",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_negedge,
	 PulseWidthHigh		=> tpw_EN_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  True, 
	 HeaderMsg		=> InstancePath & "LD",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_negedge or Pviol_EN;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT EN_ipd),D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (EN_ipd'last_event, tpd_EN_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LD_VITAL of LD is
   for VITAL_ACT
   end for;
end CFG_LD_VITAL;



 ---- CELL LDB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDB is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDB :  entity is True;
 end LDB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (SET_ipd,SET, tipd_SET);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, SET_ipd,CLR_ipd,EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_EN_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_EN_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_EN_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_EN_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_negedge,
	 TimingData		=> Tmkr_D_EN_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_negedge,
	 SetupLow		=> tsetup_D_EN_negedge_negedge,
	 HoldHigh		=> thold_D_EN_posedge_negedge,
	 HoldLow		=> thold_D_EN_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) OR (SET_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/LDB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_EN_negedge,
	 TimingData		=> Tmkr_CLR_EN_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_EN_negedge_negedge,
	 Removal		=> thold_CLR_EN_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT SET_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "LDB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_SET_EN_negedge,
	 TimingData		=> Tmkr_SET_EN_negedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_EN_negedge_negedge,
	 Removal		=> thold_SET_EN_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "LDB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_negedge,
	 PulseWidthHigh		=> tpw_EN_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT SET_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "LDB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> True,
	 HeaderMsg		=> InstancePath & "LDB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=>  TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "LDB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_negedge or Tviol_SET_EN_negedge or Pviol_SET or 
		       Pviol_CLR or Pviol_EN;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),(NOT EN_ipd),D_ipd,SET_ipd));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (SET_ipd'last_event, tpd_SET_Q, true),
		    2 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    3 => (EN_ipd'last_event, tpd_EN_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDB_VITAL of LDB is
   for VITAL_ACT
   end for;
end CFG_LDB_VITAL;



 ---- CELL LDBI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDBI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDBI :  entity is True;
 end LDBI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDBI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (SET_ipd,SET, tipd_SET);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, SET_ipd,CLR_ipd,EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_EN_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_EN_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_EN_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_EN_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QBAR_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_negedge,
	 TimingData		=> Tmkr_D_EN_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_negedge,
	 SetupLow		=> tsetup_D_EN_negedge_negedge,
	 HoldHigh		=> thold_D_EN_posedge_negedge,
	 HoldLow		=> thold_D_EN_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) OR (SET_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/LDBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_EN_negedge,
	 TimingData		=> Tmkr_CLR_EN_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_EN_negedge_negedge,
	 Removal		=> thold_CLR_EN_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT SET_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "LDBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_SET_EN_negedge,
	 TimingData		=> Tmkr_SET_EN_negedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_EN_negedge_negedge,
	 Removal		=> thold_SET_EN_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "LDBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_negedge,
	 PulseWidthHigh		=> tpw_EN_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT SET_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "LDBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> True,
	 HeaderMsg		=> InstancePath & "LDBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=>  TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "LDBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_negedge or Tviol_SET_EN_negedge or Pviol_SET or 
		       Pviol_CLR or Pviol_EN;

	VitalStateTable(
	 Result => QBAR_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),(NOT EN_ipd),D_ipd,SET_ipd));
	 QBAR_zd := Violation XOR NOT QBAR_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QBAR, true),
		     1 => (SET_ipd'last_event, tpd_SET_QBAR, true),
		    2 => (CLR_ipd'last_event, tpd_CLR_QBAR, true),
		    3 => (EN_ipd'last_event, tpd_EN_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDBI_VITAL of LDBI is
   for VITAL_ACT
   end for;
end CFG_LDBI_VITAL;



 ---- CELL LDC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDC :  entity is True;
 end LDC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_EN_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_EN_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_negedge,
	 TimingData		=> Tmkr_D_EN_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_negedge,
	 SetupLow		=> tsetup_D_EN_negedge_negedge,
	 HoldHigh		=> thold_D_EN_posedge_negedge,
	 HoldLow		=> thold_D_EN_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/LDC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_EN_negedge,
	 TimingData		=> Tmkr_CLR_EN_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_EN_negedge_negedge,
	 Removal		=> thold_CLR_EN_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  True,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "LDC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_negedge,
	 PulseWidthHigh		=> tpw_EN_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "LDC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> True,
	 HeaderMsg		=> InstancePath & "LDC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_negedge or Pviol_CLR or Pviol_EN;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),(NOT EN_ipd),D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    2 => (EN_ipd'last_event, tpd_EN_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDC_VITAL of LDC is
   for VITAL_ACT
   end for;
end CFG_LDC_VITAL;



 ---- CELL LDCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDCI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDCI :  entity is True;
 end LDCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_EN_negedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_EN_negedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QBAR_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_negedge,
	 TimingData		=> Tmkr_D_EN_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_negedge,
	 SetupLow		=> tsetup_D_EN_negedge_negedge,
	 HoldHigh		=> thold_D_EN_posedge_negedge,
	 HoldLow		=> thold_D_EN_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/LDCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_EN_negedge,
	 TimingData		=> Tmkr_CLR_EN_negedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_EN_negedge_negedge,
	 Removal		=> thold_CLR_EN_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  True,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "LDCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_negedge,
	 PulseWidthHigh		=> tpw_EN_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "LDCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> True,
	 HeaderMsg		=> InstancePath & "LDCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_negedge or Pviol_CLR or Pviol_EN;

	VitalStateTable(
	 Result => QBAR_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),(NOT EN_ipd),D_ipd,'0'));
	 QBAR_zd := Violation XOR NOT QBAR_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QBAR, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_QBAR, true),
		    2 => (EN_ipd'last_event, tpd_EN_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDCI_VITAL of LDCI is
   for VITAL_ACT
   end for;
end CFG_LDCI_VITAL;



 ---- CELL LDI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDI :  entity is True;
 end LDI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QBAR_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_negedge,
	 TimingData		=> Tmkr_D_EN_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_negedge,
	 SetupLow		=> tsetup_D_EN_negedge_negedge,
	 HoldHigh		=> thold_D_EN_posedge_negedge,
	 HoldLow		=> thold_D_EN_negedge_negedge,
	 CheckEnabled		=>  True, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/LDI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_negedge,
	 PulseWidthHigh		=> tpw_EN_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  True, 
	 HeaderMsg		=> InstancePath & "LDI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_negedge or Pviol_EN;

	VitalStateTable(
	 Result => QBAR_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT EN_ipd),D_ipd,'0'));
	 QBAR_zd := Violation XOR NOT QBAR_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QBAR, true),
		    1 => (EN_ipd'last_event, tpd_EN_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDI_VITAL of LDI is
   for VITAL_ACT
   end for;
end CFG_LDI_VITAL;



 ---- CELL LDL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDL is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDL :  entity is True;
 end LDL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_posedge,
	 TimingData		=> Tmkr_D_EN_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_posedge,
	 SetupLow		=> tsetup_D_EN_negedge_posedge,
	 HoldHigh		=> thold_D_EN_posedge_posedge,
	 HoldLow		=> thold_D_EN_negedge_posedge,
	 CheckEnabled		=>  True, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/LDL",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_EN_negedge,
	 CheckEnabled		=>  True, 
	 HeaderMsg		=> InstancePath & "LDL",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_posedge or Pviol_EN;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',EN_ipd,D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (EN_ipd'last_event, tpd_EN_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDL_VITAL of LDL is
   for VITAL_ACT
   end for;
end CFG_LDL_VITAL;



 ---- CELL LDLB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDLB is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDLB :  entity is True;
 end LDLB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDLB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (SET_ipd,SET, tipd_SET);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, SET_ipd,CLR_ipd,EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_EN_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_EN_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_EN_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_EN_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_posedge,
	 TimingData		=> Tmkr_D_EN_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_posedge,
	 SetupLow		=> tsetup_D_EN_negedge_posedge,
	 HoldHigh		=> thold_D_EN_posedge_posedge,
	 HoldLow		=> thold_D_EN_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) OR (SET_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/LDLB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_EN_posedge,
	 TimingData		=> Tmkr_CLR_EN_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_EN_negedge_posedge,
	 Removal		=> thold_CLR_EN_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT SET_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "LDLB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_SET_EN_posedge,
	 TimingData		=> Tmkr_SET_EN_posedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_EN_negedge_posedge,
	 Removal		=> thold_SET_EN_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "LDLB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_EN_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT SET_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "LDLB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> True,
	 HeaderMsg		=> InstancePath & "LDLB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=>  TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "LDLB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_posedge or Tviol_SET_EN_posedge or Pviol_SET or 
		       Pviol_CLR or Pviol_EN;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),EN_ipd,D_ipd,SET_ipd));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (SET_ipd'last_event, tpd_SET_Q, true),
		    2 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    3 => (EN_ipd'last_event, tpd_EN_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDLB_VITAL of LDLB is
   for VITAL_ACT
   end for;
end CFG_LDLB_VITAL;



 ---- CELL LDLBI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDLBI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDLBI :  entity is True;
 end LDLBI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDLBI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (SET_ipd,SET, tipd_SET);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, SET_ipd,CLR_ipd,EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_EN_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_EN_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_EN_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_EN_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QBAR_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_posedge,
	 TimingData		=> Tmkr_D_EN_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_posedge,
	 SetupLow		=> tsetup_D_EN_negedge_posedge,
	 HoldHigh		=> thold_D_EN_posedge_posedge,
	 HoldLow		=> thold_D_EN_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) OR (SET_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/LDLBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_EN_posedge,
	 TimingData		=> Tmkr_CLR_EN_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_EN_negedge_posedge,
	 Removal		=> thold_CLR_EN_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT SET_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "LDLBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_SET_EN_posedge,
	 TimingData		=> Tmkr_SET_EN_posedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_EN_negedge_posedge,
	 Removal		=> thold_SET_EN_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "LDLBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_EN_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT SET_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "LDLBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> True,
	 HeaderMsg		=> InstancePath & "LDLBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=>  TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "LDLBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_posedge or Tviol_SET_EN_posedge or Pviol_SET or 
		       Pviol_CLR or Pviol_EN;

	VitalStateTable(
	 Result => QBAR_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),EN_ipd,D_ipd,SET_ipd));
	 QBAR_zd := Violation XOR NOT QBAR_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QBAR, true),
		     1 => (SET_ipd'last_event, tpd_SET_QBAR, true),
		    2 => (CLR_ipd'last_event, tpd_CLR_QBAR, true),
		    3 => (EN_ipd'last_event, tpd_EN_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDLBI_VITAL of LDLBI is
   for VITAL_ACT
   end for;
end CFG_LDLBI_VITAL;



 ---- CELL LDLC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDLC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDLC :  entity is True;
 end LDLC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDLC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_EN_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_EN_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_posedge,
	 TimingData		=> Tmkr_D_EN_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_posedge,
	 SetupLow		=> tsetup_D_EN_negedge_posedge,
	 HoldHigh		=> thold_D_EN_posedge_posedge,
	 HoldLow		=> thold_D_EN_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/LDLC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_EN_posedge,
	 TimingData		=> Tmkr_CLR_EN_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_EN_negedge_posedge,
	 Removal		=> thold_CLR_EN_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  True,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "LDLC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_EN_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "LDLC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> True,
	 HeaderMsg		=> InstancePath & "LDLC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_posedge or Pviol_CLR or Pviol_EN;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),EN_ipd,D_ipd,'0'));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_Q, true),
		    2 => (EN_ipd'last_event, tpd_EN_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDLC_VITAL of LDLC is
   for VITAL_ACT
   end for;
end CFG_LDLC_VITAL;



 ---- CELL LDLCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDLCI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		CLR		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDLCI :  entity is True;
 end LDLCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDLCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, CLR_ipd,EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_EN_posedge	: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_EN_posedge         : VitalTimingDataType	:= VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QBAR_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_posedge,
	 TimingData		=> Tmkr_D_EN_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_posedge,
	 SetupLow		=> tsetup_D_EN_negedge_posedge,
	 HoldHigh		=> thold_D_EN_posedge_posedge,
	 HoldLow		=> thold_D_EN_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((CLR_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/LDLCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_CLR_EN_posedge,
	 TimingData		=> Tmkr_CLR_EN_posedge,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_CLR_EN_negedge_posedge,
	 Removal		=> thold_CLR_EN_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  True,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "LDLCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_EN_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "LDLCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData		=> PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> True,
	 HeaderMsg		=> InstancePath & "LDLCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_posedge or Pviol_CLR or Pviol_EN;

	VitalStateTable(
	 Result => QBAR_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		 (NOT CLR_ipd),EN_ipd,D_ipd,'0'));
	 QBAR_zd := Violation XOR NOT QBAR_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QBAR, true),
		    1 => (CLR_ipd'last_event, tpd_CLR_QBAR, true),
		    2 => (EN_ipd'last_event, tpd_EN_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDLCI_VITAL of LDLCI is
   for VITAL_ACT
   end for;
end CFG_LDLCI_VITAL;



 ---- CELL LDLI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDLI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDLI :  entity is True;
 end LDLI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDLI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QBAR_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_posedge,
	 TimingData		=> Tmkr_D_EN_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_posedge,
	 SetupLow		=> tsetup_D_EN_negedge_posedge,
	 HoldHigh		=> thold_D_EN_posedge_posedge,
	 HoldLow		=> thold_D_EN_negedge_posedge,
	 CheckEnabled		=>  True, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/LDLI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_EN_negedge,
	 CheckEnabled		=>  True, 
	 HeaderMsg		=> InstancePath & "LDLI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_posedge or Pviol_EN;

	VitalStateTable(
	 Result => QBAR_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',EN_ipd,D_ipd,'0'));
	 QBAR_zd := Violation XOR NOT QBAR_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QBAR, true),
		    1 => (EN_ipd'last_event, tpd_EN_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDLI_VITAL of LDLI is
   for VITAL_ACT
   end for;
end CFG_LDLI_VITAL;



 ---- CELL LDLS ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDLS is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDLS :  entity is True;
 end LDLS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDLS is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (SET_ipd,SET, tipd_SET);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, SET_ipd,EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_EN_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_EN_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_posedge,
	 TimingData		=> Tmkr_D_EN_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_posedge,
	 SetupLow		=> tsetup_D_EN_negedge_posedge,
	 HoldHigh		=> thold_D_EN_posedge_posedge,
	 HoldLow		=> thold_D_EN_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((SET_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/LDLS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_SET_EN_posedge,
	 TimingData		=> Tmkr_SET_EN_posedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_EN_negedge_posedge,
	 Removal		=> thold_SET_EN_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  True,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "LDLS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_EN_negedge,
	 CheckEnabled		=>  TO_X01(((NOT SET_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "LDLS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 	True,
	 HeaderMsg		=> InstancePath & "LDLS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_posedge or Tviol_SET_EN_posedge or Pviol_SET or 
		       Pviol_EN;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',EN_ipd,D_ipd,SET_ipd));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (SET_ipd'last_event, tpd_SET_Q, true),
		    2 => (EN_ipd'last_event, tpd_EN_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDLS_VITAL of LDLS is
   for VITAL_ACT
   end for;
end CFG_LDLS_VITAL;



 ---- CELL LDLSI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDLSI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_posedge		:  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_negedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDLSI :  entity is True;
 end LDLSI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDLSI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (SET_ipd,SET, tipd_SET);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, SET_ipd,EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_EN_posedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_EN_posedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QBAR_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_posedge,
	 TimingData		=> Tmkr_D_EN_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_posedge,
	 SetupLow		=> tsetup_D_EN_negedge_posedge,
	 HoldHigh		=> thold_D_EN_posedge_posedge,
	 HoldLow		=> thold_D_EN_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((SET_ipd) ) ) /= '1', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/LDLSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_SET_EN_posedge,
	 TimingData		=> Tmkr_SET_EN_posedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_EN_negedge_posedge,
	 Removal		=> thold_SET_EN_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  True,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "LDLSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_posedge,
	 PulseWidthHigh         => 0 ns,
	 PulseWidthLow		=> tpw_EN_negedge,
	 CheckEnabled		=>  TO_X01(((NOT SET_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "LDLSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 	True,
	 HeaderMsg		=> InstancePath & "LDLSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_posedge or Tviol_SET_EN_posedge or Pviol_SET or 
		       Pviol_EN;

	VitalStateTable(
	 Result => QBAR_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',EN_ipd,D_ipd,SET_ipd));
	 QBAR_zd := Violation XOR NOT QBAR_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QBAR, true),
		     1 => (SET_ipd'last_event, tpd_SET_QBAR, true),
		    2 => (EN_ipd'last_event, tpd_EN_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDLSI_VITAL of LDLSI is
   for VITAL_ACT
   end for;
end CFG_LDLSI_VITAL;



 ---- CELL LDS ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDS is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDS :  entity is True;
 end LDS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDS is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (SET_ipd,SET, tipd_SET);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, SET_ipd,EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_EN_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_EN_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS Q_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_negedge,
	 TimingData		=> Tmkr_D_EN_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_negedge,
	 SetupLow		=> tsetup_D_EN_negedge_negedge,
	 HoldHigh		=> thold_D_EN_posedge_negedge,
	 HoldLow		=> thold_D_EN_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((SET_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/LDS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_SET_EN_negedge,
	 TimingData		=> Tmkr_SET_EN_negedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_EN_negedge_negedge,
	 Removal		=> thold_SET_EN_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  True,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "LDS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_negedge,
	 PulseWidthHigh		=> tpw_EN_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT SET_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "LDS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 	True,
	 HeaderMsg		=> InstancePath & "LDS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_negedge or Tviol_SET_EN_negedge or Pviol_SET or 
		       Pviol_EN;

	VitalStateTable(
	 Result => Q_zd,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT EN_ipd),D_ipd,SET_ipd));
	 Q_zd := Violation XOR Q_zd;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_Q, true),
		     1 => (SET_ipd'last_event, tpd_SET_Q, true),
		    2 => (EN_ipd'last_event, tpd_EN_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDS_VITAL of LDS is
   for VITAL_ACT
   end for;
end CFG_LDS_VITAL;



 ---- CELL LDSI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity LDSI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_D_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_EN_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tperiod_EN_negedge		:VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_EN_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns));


     port(
		D		:  in    STD_ULOGIC;
		SET		:  in    STD_ULOGIC;
		EN		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of LDSI :  entity is True;
 end LDSI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of LDSI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (D_ipd, D, tipd_D);
	VitalWireDelay (SET_ipd,SET, tipd_SET);
	VitalWireDelay (EN_ipd,EN, tipd_EN);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
	VITALBehavior : process (D_ipd, SET_ipd,EN_ipd)

	-- timing check results
	VARIABLE Tviol_D_EN_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_D_EN_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_EN_negedge         : STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_EN_negedge         : VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_EN	: STD_ULOGIC := '0';
	VARIABLE PInfo_EN	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q	: STD_LOGIC_VECTOR(0 to 3);
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)	:= (others => 'X');
	ALIAS QBAR_zd	:  STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData	: VitalGlitchDataType;

	begin

	------------------------
	--  Timing Check Section
	------------------------
	if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_EN_negedge,
	 TimingData		=> Tmkr_D_EN_negedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_EN_posedge_negedge,
	 SetupLow		=> tsetup_D_EN_negedge_negedge,
	 HoldHigh		=> thold_D_EN_posedge_negedge,
	 HoldLow		=> thold_D_EN_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((SET_ipd) ) ) /= '1', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/LDSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation		=> Tviol_SET_EN_negedge,
	 TimingData		=> Tmkr_SET_EN_negedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> EN_ipd,
	 RefSignalName		=> "EN",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_EN_negedge_negedge,
	 Removal		=> thold_SET_EN_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled		=>  True,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "LDSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_EN,
	 PeriodData		=> PInfo_EN,
	 TestSignal		=> EN_ipd,
	 TestSignalName		=> "EN",
	 TestDelay		=> 0 ns,
	 Period		 => tperiod_EN_negedge,
	 PulseWidthHigh		=> tpw_EN_posedge,
	 PulseWidthLow          => 0 ns,
	 CheckEnabled		=>  TO_X01(((NOT SET_ipd) ) ) /= '0', 
	 HeaderMsg		=> InstancePath & "LDSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		        => 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 	True,
	 HeaderMsg		=> InstancePath & "LDSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

   end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_EN_negedge or Tviol_SET_EN_negedge or Pviol_SET or 
		       Pviol_EN;

	VitalStateTable(
	 Result => QBAR_temp,
	 PreviousDataIn => PrevData_Q,
	 StateTable => dlatch_DL2C_Q_tab,
	 DataIn => (
		'1',(NOT EN_ipd),D_ipd,SET_ipd));
	 QBAR_zd := Violation XOR NOT QBAR_temp;
	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (D_ipd'last_event, tpd_D_QBAR, true),
		     1 => (SET_ipd'last_event, tpd_SET_QBAR, true),
		    2 => (EN_ipd'last_event, tpd_EN_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_LDSI_VITAL of LDSI is
   for VITAL_ACT
   end for;
end CFG_LDSI_VITAL;



 ---- CELL MUX2H ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MUX2H is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MUX2H :  entity is True;
 end MUX2H;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of MUX2H is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( A_ipd , B_ipd , (NOT S_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (S_ipd'last_event,tpd_S_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MUX2H_VITAL of MUX2H is 
    for VITAL_ACT
    end for;
 end CFG_MUX2H_VITAL;



 ---- CELL MUX2L ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity MUX2L is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_S_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_S		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		S		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of MUX2L :  entity is True;
 end MUX2L;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of MUX2L is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL S_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (S_ipd, S, tipd_S);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, S_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( A_ipd , B_ipd , S_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (S_ipd'last_event,tpd_S_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_MUX2L_VITAL of MUX2L is 
    for VITAL_ACT
    end for;
 end CFG_MUX2L_VITAL;



 ---- CELL NAND2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND2 :  entity is True;
 end NAND2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of NAND2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT A_ipd)  OR  (NOT B_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND2_VITAL of NAND2 is 
    for VITAL_ACT
    end for;
 end CFG_NAND2_VITAL;



 ---- CELL NAND2FT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND2FT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND2FT :  entity is True;
 end NAND2FT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of NAND2FT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( A_ipd  OR  (NOT B_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND2FT_VITAL of NAND2FT is 
    for VITAL_ACT
    end for;
 end CFG_NAND2FT_VITAL;



 ---- CELL NAND3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND3 :  entity is True;
 end NAND3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of NAND3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND3_VITAL of NAND3 is 
    for VITAL_ACT
    end for;
 end CFG_NAND3_VITAL;



 ---- CELL NAND3FFT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND3FFT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND3FFT :  entity is True;
 end NAND3FFT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of NAND3FFT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  OR  B_ipd ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND3FFT_VITAL of NAND3FFT is 
    for VITAL_ACT
    end for;
 end CFG_NAND3FFT_VITAL;



 ---- CELL NAND3FTT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NAND3FTT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NAND3FTT :  entity is True;
 end NAND3FTT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of NAND3FTT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  OR  (NOT B_ipd) ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NAND3FTT_VITAL of NAND3FTT is 
    for VITAL_ACT
    end for;
 end CFG_NAND3FTT_VITAL;



 ---- CELL NOR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR2 :  entity is True;
 end NOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of NOR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT A_ipd)  AND  (NOT B_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR2_VITAL of NOR2 is 
    for VITAL_ACT
    end for;
 end CFG_NOR2_VITAL;



 ---- CELL NOR2FT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR2FT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR2FT :  entity is True;
 end NOR2FT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of NOR2FT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( A_ipd  AND  (NOT B_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR2FT_VITAL of NOR2FT is 
    for VITAL_ACT
    end for;
 end CFG_NOR2FT_VITAL;



 ---- CELL NOR3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR3 :  entity is True;
 end NOR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of NOR3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT B_ipd) ) AND  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR3_VITAL of NOR3 is 
    for VITAL_ACT
    end for;
 end CFG_NOR3_VITAL;



 ---- CELL NOR3FFT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR3FFT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR3FFT :  entity is True;
 end NOR3FFT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of NOR3FFT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  B_ipd ) AND  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR3FFT_VITAL of NOR3FFT is 
    for VITAL_ACT
    end for;
 end CFG_NOR3FFT_VITAL;



 ---- CELL NOR3FTT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NOR3FTT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NOR3FTT :  entity is True;
 end NOR3FTT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of NOR3FTT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  (NOT B_ipd) ) AND  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NOR3FTT_VITAL of NOR3FTT is 
    for VITAL_ACT
    end for;
 end CFG_NOR3FTT_VITAL;



 ---- CELL NUBBLE ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity NUBBLE is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of NUBBLE :  entity is True;
 end NUBBLE;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of NUBBLE is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_NUBBLE_VITAL of NUBBLE is 
    for VITAL_ACT
    end for;
 end CFG_NUBBLE_VITAL;



 ---- CELL OA21 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA21 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA21 :  entity is True;
 end OA21;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OA21 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, C_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  C_ipd ) OR ( B_ipd  AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (C_ipd'last_event,tpd_C_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA21_VITAL of OA21 is 
    for VITAL_ACT
    end for;
 end CFG_OA21_VITAL;



 ---- CELL OA21FTF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA21FTF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA21FTF :  entity is True;
 end OA21FTF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OA21FTF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, C_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT C_ipd) ) OR ( B_ipd  AND  (NOT C_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (C_ipd'last_event,tpd_C_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA21FTF_VITAL of OA21FTF is 
    for VITAL_ACT
    end for;
 end CFG_OA21FTF_VITAL;



 ---- CELL OA21FTT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA21FTT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA21FTT :  entity is True;
 end OA21FTT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OA21FTT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, C_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  C_ipd ) OR ( B_ipd  AND  C_ipd ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (C_ipd'last_event,tpd_C_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA21FTT_VITAL of OA21FTT is 
    for VITAL_ACT
    end for;
 end CFG_OA21FTT_VITAL;



 ---- CELL OA21TTF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OA21TTF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OA21TTF :  entity is True;
 end OA21TTF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OA21TTF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, C_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  (NOT C_ipd) ) OR ( B_ipd  AND  (NOT C_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (C_ipd'last_event,tpd_C_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OA21TTF_VITAL of OA21TTF is 
    for VITAL_ACT
    end for;
 end CFG_OA21TTF_VITAL;



 ---- CELL OAI21 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OAI21 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OAI21 :  entity is True;
 end OAI21;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OAI21 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  AND  (NOT B_ipd) ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OAI21_VITAL of OAI21 is 
    for VITAL_ACT
    end for;
 end CFG_OAI21_VITAL;



 ---- CELL OAI21FTF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OAI21FTF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OAI21FTF :  entity is True;
 end OAI21FTF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OAI21FTF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  (NOT B_ipd) ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OAI21FTF_VITAL of OAI21FTF is 
    for VITAL_ACT
    end for;
 end CFG_OAI21FTF_VITAL;



 ---- CELL OAI21FTT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OAI21FTT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OAI21FTT :  entity is True;
 end OAI21FTT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OAI21FTT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  AND  (NOT B_ipd) ) OR  (NOT C_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OAI21FTT_VITAL of OAI21FTT is 
    for VITAL_ACT
    end for;
 end CFG_OAI21FTT_VITAL;



 ---- CELL OAI21TTF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OAI21TTF is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		C		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OAI21TTF :  entity is True;
 end OAI21TTF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OAI21TTF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL C_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (C_ipd, C, tipd_C);
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (C_ipd, A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( C_ipd  OR ( (NOT A_ipd)  AND  (NOT B_ipd) ));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (C_ipd'last_event,tpd_C_Y, true),
	             1 => (A_ipd'last_event,tpd_A_Y, true),
	             2 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OAI21TTF_VITAL of OAI21TTF is 
    for VITAL_ACT
    end for;
 end CFG_OAI21TTF_VITAL;



 ---- CELL OB25HH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB25HH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB25HH :  entity is True;
 end OB25HH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB25HH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB25HH_VITAL of OB25HH is 
    for VITAL_ACT
    end for;
 end CFG_OB25HH_VITAL;



 ---- CELL OB25HL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB25HL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB25HL :  entity is True;
 end OB25HL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB25HL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB25HL_VITAL of OB25HL is 
    for VITAL_ACT
    end for;
 end CFG_OB25HL_VITAL;



 ---- CELL OB25HN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB25HN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB25HN :  entity is True;
 end OB25HN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB25HN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB25HN_VITAL of OB25HN is 
    for VITAL_ACT
    end for;
 end CFG_OB25HN_VITAL;



 ---- CELL OB25LH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB25LH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB25LH :  entity is True;
 end OB25LH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB25LH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB25LH_VITAL of OB25LH is 
    for VITAL_ACT
    end for;
 end CFG_OB25LH_VITAL;



 ---- CELL OB25LL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB25LL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB25LL :  entity is True;
 end OB25LL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB25LL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB25LL_VITAL of OB25LL is 
    for VITAL_ACT
    end for;
 end CFG_OB25LL_VITAL;



 ---- CELL OB25LN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB25LN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB25LN :  entity is True;
 end OB25LN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB25LN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB25LN_VITAL of OB25LN is 
    for VITAL_ACT
    end for;
 end CFG_OB25LN_VITAL;



 ---- CELL OB25LPHH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB25LPHH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB25LPHH :  entity is True;
 end OB25LPHH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB25LPHH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB25LPHH_VITAL of OB25LPHH is 
    for VITAL_ACT
    end for;
 end CFG_OB25LPHH_VITAL;



 ---- CELL OB25LPHL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB25LPHL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB25LPHL :  entity is True;
 end OB25LPHL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB25LPHL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB25LPHL_VITAL of OB25LPHL is 
    for VITAL_ACT
    end for;
 end CFG_OB25LPHL_VITAL;



 ---- CELL OB25LPHN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB25LPHN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB25LPHN :  entity is True;
 end OB25LPHN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB25LPHN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB25LPHN_VITAL of OB25LPHN is 
    for VITAL_ACT
    end for;
 end CFG_OB25LPHN_VITAL;



 ---- CELL OB25LPLH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB25LPLH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB25LPLH :  entity is True;
 end OB25LPLH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB25LPLH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB25LPLH_VITAL of OB25LPLH is 
    for VITAL_ACT
    end for;
 end CFG_OB25LPLH_VITAL;



 ---- CELL OB25LPLL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB25LPLL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB25LPLL :  entity is True;
 end OB25LPLL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB25LPLL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB25LPLL_VITAL of OB25LPLL is 
    for VITAL_ACT
    end for;
 end CFG_OB25LPLL_VITAL;



 ---- CELL OB25LPLN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB25LPLN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB25LPLN :  entity is True;
 end OB25LPLN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB25LPLN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB25LPLN_VITAL of OB25LPLN is 
    for VITAL_ACT
    end for;
 end CFG_OB25LPLN_VITAL;



 ---- CELL OB33LH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB33LH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB33LH :  entity is True;
 end OB33LH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB33LH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB33LH_VITAL of OB33LH is 
    for VITAL_ACT
    end for;
 end CFG_OB33LH_VITAL;



 ---- CELL OB33LL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB33LL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB33LL :  entity is True;
 end OB33LL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB33LL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB33LL_VITAL of OB33LL is 
    for VITAL_ACT
    end for;
 end CFG_OB33LL_VITAL;



 ---- CELL OB33LN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB33LN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB33LN :  entity is True;
 end OB33LN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB33LN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB33LN_VITAL of OB33LN is 
    for VITAL_ACT
    end for;
 end CFG_OB33LN_VITAL;



 ---- CELL OB33PH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB33PH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB33PH :  entity is True;
 end OB33PH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB33PH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB33PH_VITAL of OB33PH is 
    for VITAL_ACT
    end for;
 end CFG_OB33PH_VITAL;



 ---- CELL OB33PL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB33PL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB33PL :  entity is True;
 end OB33PL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB33PL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB33PL_VITAL of OB33PL is 
    for VITAL_ACT
    end for;
 end CFG_OB33PL_VITAL;



 ---- CELL OB33PN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OB33PN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OB33PN :  entity is True;
 end OB33PN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OB33PN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OB33PN_VITAL of OB33PN is 
    for VITAL_ACT
    end for;
 end CFG_OB33PN_VITAL;



 ---- CELL OR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR2 :  entity is True;
 end OR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( A_ipd  OR  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR2_VITAL of OR2 is 
    for VITAL_ACT
    end for;
 end CFG_OR2_VITAL;



 ---- CELL OR2FT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR2FT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR2FT :  entity is True;
 end OR2FT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OR2FT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := ( (NOT A_ipd)  OR  B_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR2FT_VITAL of OR2FT is 
    for VITAL_ACT
    end for;
 end CFG_OR2FT_VITAL;



 ---- CELL OR3 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR3 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR3 :  entity is True;
 end OR3;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OR3 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( A_ipd  OR  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR3_VITAL of OR3 is 
    for VITAL_ACT
    end for;
 end CFG_OR3_VITAL;



 ---- CELL OR3FFT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR3FFT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR3FFT :  entity is True;
 end OR3FFT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OR3FFT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  OR  (NOT B_ipd) ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR3FFT_VITAL of OR3FFT is 
    for VITAL_ACT
    end for;
 end CFG_OR3FFT_VITAL;



 ---- CELL OR3FTT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OR3FTT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_C_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_C		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		C		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OR3FTT :  entity is True;
 end OR3FTT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OR3FTT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';
	SIGNAL C_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	VitalWireDelay (C_ipd, C, tipd_C);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd, C_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd := (( (NOT A_ipd)  OR  B_ipd ) OR  C_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true),
	             2 => (C_ipd'last_event,tpd_C_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_OR3FTT_VITAL of OR3FTT is 
    for VITAL_ACT
    end for;
 end CFG_OR3FTT_VITAL;



 ---- CELL PWR ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity PWR is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True		);
    port(
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of PWR :  entity is True;
 end PWR;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of PWR is
	attribute VITAL_LEVEL0 of VITAL_ACT : architecture is True;


begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	--- Empty
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
        Y<= '1';


end VITAL_ACT;

 configuration CFG_PWR_VITAL of PWR is 
    for VITAL_ACT
    end for;
 end CFG_PWR_VITAL;



 ---- CELL XNOR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XNOR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XNOR2 :  entity is True;
 end XNOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of XNOR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XNOR2_VITAL of XNOR2 is 
    for VITAL_ACT
    end for;
 end CFG_XNOR2_VITAL;



 ---- CELL XNOR2FT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XNOR2FT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XNOR2FT :  entity is True;
 end XNOR2FT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of XNOR2FT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  NOT VitalMUX2( B_ipd , (NOT B_ipd) , A_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XNOR2FT_VITAL of XNOR2FT is 
    for VITAL_ACT
    end for;
 end CFG_XNOR2FT_VITAL;



 ---- CELL XOR2 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XOR2 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XOR2 :  entity is True;
 end XOR2;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of XOR2 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( B_ipd , (NOT B_ipd) , (NOT A_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XOR2_VITAL of XOR2 is 
    for VITAL_ACT
    end for;
 end CFG_XOR2_VITAL;



 ---- CELL XOR2FT ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity XOR2FT is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_B_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_B		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		B		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of XOR2FT :  entity is True;
 end XOR2FT;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of XOR2FT is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL B_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (B_ipd, B, tipd_B);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, B_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       Y_zd :=  VitalMUX2( B_ipd , (NOT B_ipd) , A_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (B_ipd'last_event,tpd_B_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_XOR2FT_VITAL of XOR2FT is 
    for VITAL_ACT
    end for;
 end CFG_XOR2FT_VITAL;



 ---- CELL DFF ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFF is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFF :  entity is True;
 end DFF;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFF is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  True, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFF",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>True,
	 HeaderMsg		=> InstancePath & "DFF",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, '0', '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFF_VITAL of DFF is
   for VITAL_ACT
   end for;
end CFG_DFF_VITAL;



 ---- CELL DFFB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFB is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFB :  entity is True;
 end DFFB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (SET_ipd,SET, tipd_SET);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, SET_ipd,CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT SET_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFFB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_SET_CLK_posedge,
	 TimingData		=> Tmkr_SET_CLK_posedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_CLK_negedge_posedge,
	 Removal		=> thold_SET_CLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFFB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_posedge,
	 Removal               => thold_CLR_CLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01(( NOT SET_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFFB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((NOT SET_ipd) AND ( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFFB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => True,
	 HeaderMsg              => InstancePath & "DFFB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 		TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFFB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_SET_CLK_posedge or 
	 Tviol_SET_CLK_posedge or Pviol_SET or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_delayed, Q_zd, D_delayed, '0', (NOT SET_ipd), CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (SET_ipd'last_event, tpd_SET_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFB_VITAL of DFFB is
   for VITAL_ACT
   end for;
end CFG_DFFB_VITAL;



 ---- CELL DFFBI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFBI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFBI :  entity is True;
 end DFFBI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFBI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (SET_ipd,SET, tipd_SET);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, SET_ipd,CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QBAR_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT SET_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFFBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_SET_CLK_posedge,
	 TimingData		=> Tmkr_SET_CLK_posedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_CLK_negedge_posedge,
	 Removal		=> thold_SET_CLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFFBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_posedge,
	 Removal               => thold_CLR_CLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01(( NOT SET_ipd)) /= '0',
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFFBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((NOT SET_ipd) AND ( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFFBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => True,
	 HeaderMsg              => InstancePath & "DFFBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 		TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFFBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_SET_CLK_posedge or 
	 Tviol_SET_CLK_posedge or Pviol_SET or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => QBAR_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_delayed, QBAR_temp, D_delayed, '0', (NOT SET_ipd), CLK_ipd));
   QBAR_zd := Violation XOR  (NOT QBAR_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QBAR, true),
	             1=> (SET_ipd'last_event, tpd_SET_QBAR, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFBI_VITAL of DFFBI is
   for VITAL_ACT
   end for;
end CFG_DFFBI_VITAL;



 ---- CELL DFFC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFC :  entity is True;
 end DFFC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFFC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_posedge,
	 Removal               => thold_CLR_CLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>    True,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFFC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFFC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => True,
	 HeaderMsg              => InstancePath & "DFFC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_delayed, Q_zd, D_delayed, '0', '1', CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFC_VITAL of DFFC is
   for VITAL_ACT
   end for;
end CFG_DFFC_VITAL;



 ---- CELL DFFCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFCI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFCI :  entity is True;
 end DFFCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QBAR_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFFCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_posedge,
	 TimingData             => Tmkr_CLR_CLK_posedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_posedge,
	 Removal               => thold_CLR_CLK_negedge_posedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>    True,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFFCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFFCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => True,
	 HeaderMsg              => InstancePath & "DFFCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QBAR_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_delayed, QBAR_temp, D_delayed, '0', '1', CLK_ipd));
   QBAR_zd := Violation XOR  (NOT QBAR_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QBAR, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFCI_VITAL of DFFCI is
   for VITAL_ACT
   end for;
end CFG_DFFCI_VITAL;



 ---- CELL DFFI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFI :  entity is True;
 end DFFI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QBAR_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  True, 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFFI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>True,
	 HeaderMsg		=> InstancePath & "DFFI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QBAR_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, QBAR_temp, D_delayed, '0', '1', CLK_ipd));
   QBAR_zd := Violation XOR  (NOT QBAR_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFI_VITAL of DFFI is
   for VITAL_ACT
   end for;
end CFG_DFFI_VITAL;



 ---- CELL DFFL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFL is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFL :  entity is True;
 end DFFL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  True, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFFL",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>True,
	 HeaderMsg		=> InstancePath & "DFFL",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed, '0', '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFL_VITAL of DFFL is
   for VITAL_ACT
   end for;
end CFG_DFFL_VITAL;



 ---- CELL DFFLB ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFLB is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFLB :  entity is True;
 end DFFLB;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFLB is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (SET_ipd,SET, tipd_SET);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, SET_ipd,CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT SET_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFFLB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_SET_CLK_negedge,
	 TimingData		=> Tmkr_SET_CLK_negedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_CLK_negedge_negedge,
	 Removal		=> thold_SET_CLK_negedge_negedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFFLB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_negedge,
	 Removal               => thold_CLR_CLK_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01(( NOT SET_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFFLB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT SET_ipd) AND ( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFFLB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => True,
	 HeaderMsg              => InstancePath & "DFFLB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 		TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFFLB",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_SET_CLK_negedge or 
	 Tviol_SET_CLK_negedge or Pviol_SET or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_ipd, Q_zd, D_delayed, '0', (NOT SET_ipd), CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (SET_ipd'last_event, tpd_SET_Q, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFLB_VITAL of DFFLB is
   for VITAL_ACT
   end for;
end CFG_DFFLB_VITAL;



 ---- CELL DFFLBI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFLBI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFLBI :  entity is True;
 end DFFLBI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFLBI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (SET_ipd,SET, tipd_SET);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, SET_ipd,CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QBAR_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) AND (NOT SET_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFFLBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_SET_CLK_negedge,
	 TimingData		=> Tmkr_SET_CLK_negedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_CLK_negedge_negedge,
	 Removal		=> thold_SET_CLK_negedge_negedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  TO_X01(( NOT CLR_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFFLBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_negedge,
	 Removal               => thold_CLR_CLK_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>      TO_X01(( NOT SET_ipd)) /= '0',
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFFLBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT SET_ipd) AND ( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFFLBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => True,
	 HeaderMsg              => InstancePath & "DFFLBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 		TO_X01( NOT CLR_ipd) /='0',
	 HeaderMsg		=> InstancePath & "DFFLBI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_SET_CLK_negedge or 
	 Tviol_SET_CLK_negedge or Pviol_SET or Pviol_CLR or Pviol_CLK;

  VitalStateTable(
   Result => QBAR_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_ipd, QBAR_temp, D_delayed, '0', (NOT SET_ipd), CLK_delayed));
   QBAR_zd := Violation XOR  (NOT QBAR_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QBAR, true),
	             1=> (SET_ipd'last_event, tpd_SET_QBAR, true),
	            2=> (CLR_ipd'last_event, tpd_CLR_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFLBI_VITAL of DFFLBI is
   for VITAL_ACT
   end for;
end CFG_DFFLBI_VITAL;



 ---- CELL DFFLC ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFLC is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFLC :  entity is True;
 end DFFLC;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFLC is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFFLC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_negedge,
	 Removal               => thold_CLR_CLK_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>    True,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFFLC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFFLC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => True,
	 HeaderMsg              => InstancePath & "DFFLC",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_ipd, Q_zd, D_delayed, '0', '1', CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFLC_VITAL of DFFLC is
   for VITAL_ACT
   end for;
end CFG_DFFLC_VITAL;



 ---- CELL DFFLCI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFLCI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLR_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_CLR_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_CLR_posedge		:  VitalDelayType := 0.000 ns;
		tipd_CLR		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLR		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFLCI :  entity is True;
 end DFFLCI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFLCI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLR_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLR_ipd,CLR, tipd_CLR);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLR_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_CLR_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_CLR_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_CLR	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLR	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QBAR_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT CLR_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFFLCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck (
	 Violation              => Tviol_CLR_CLK_negedge,
	 TimingData             => Tmkr_CLR_CLK_negedge,
	 TestSignal             => CLR_ipd,
	 TestSignalName         => "CLR",
	 TestDelay              => 0 ns,
	 RefSignal              => CLK_ipd,
	 RefSignalName          => "CLK",
	 RefDelay               => 0 ns,
	 Recovery              => trecovery_CLR_CLK_negedge_negedge,
	 Removal               => thold_CLR_CLK_negedge_negedge,
	 ActiveLow		=> FALSE,
	 CheckEnabled           =>    True,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFFLCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01((( NOT CLR_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFFLCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLR,
	 PeriodData             => PInfo_CLR,
	 TestSignal		=> CLR_ipd,
	 TestSignalName		=> "CLR",
	 TestDelay		=> 0 ns,
	 Period			=> 0 ns,
	 PulseWidthHigh		=> tpw_CLR_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled           => True,
	 HeaderMsg              => InstancePath & "DFFLCI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLR or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QBAR_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             (NOT CLR_ipd), CLK_ipd, QBAR_temp, D_delayed, '0', '1', CLK_delayed));
   QBAR_zd := Violation XOR  (NOT QBAR_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QBAR, true),
	            1=> (CLR_ipd'last_event, tpd_CLR_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFLCI_VITAL of DFFLCI is
   for VITAL_ACT
   end for;
end CFG_DFFLCI_VITAL;



 ---- CELL DFFLI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFLI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFLI :  entity is True;
 end DFFLI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFLI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QBAR_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  True, 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFFLI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>True,
	 HeaderMsg		=> InstancePath & "DFFLI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Pviol_CLK;

  VitalStateTable(
   Result => QBAR_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, QBAR_temp, D_delayed, '0', '1', CLK_delayed));
   QBAR_zd := Violation XOR  (NOT QBAR_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFLI_VITAL of DFFLI is
   for VITAL_ACT
   end for;
end CFG_DFFLI_VITAL;



 ---- CELL DFFLS ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFLS is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFLS :  entity is True;
 end DFFLS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFLS is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (SET_ipd,SET, tipd_SET);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, SET_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT SET_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFFLS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_SET_CLK_negedge,
	 TimingData		=> Tmkr_SET_CLK_negedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_CLK_negedge_negedge,
	 Removal		=> thold_SET_CLK_negedge_negedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  True,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFFLS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT SET_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFFLS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         True,
	 HeaderMsg		=> InstancePath & "DFFLS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_SET_CLK_negedge or 
	 Tviol_SET_CLK_negedge or Pviol_SET or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, Q_zd, D_delayed, '0', (NOT SET_ipd), CLK_delayed));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (SET_ipd'last_event, tpd_SET_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFLS_VITAL of DFFLS is
   for VITAL_ACT
   end for;
end CFG_DFFLS_VITAL;



 ---- CELL DFFLSI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFLSI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_negedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_negedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFLSI :  entity is True;
 end DFFLSI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFLSI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (SET_ipd,SET, tipd_SET);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, SET_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_CLK_negedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_CLK_negedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QBAR_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_negedge, 
	 TimingData		=> Tmkr_D_CLK_negedge, 
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_negedge,
	 SetupLow		=> tsetup_D_CLK_negedge_negedge,
	 HoldHigh		=> thold_D_CLK_posedge_negedge,
	 HoldLow		=> thold_D_CLK_negedge_negedge,
	 CheckEnabled		=>  TO_X01(((NOT SET_ipd) ) ) /= '0', 
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "/DFFLSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_SET_CLK_negedge,
	 TimingData		=> Tmkr_SET_CLK_negedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_CLK_negedge_negedge,
	 Removal		=> thold_SET_CLK_negedge_negedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  True,
	 RefTransition		=> 'F',
	 HeaderMsg		=> InstancePath & "DFFLSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_negedge,
	 CheckEnabled		=>		TO_X01(((NOT SET_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFFLSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         True,
	 HeaderMsg		=> InstancePath & "DFFLSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_negedge or 
	 Tviol_SET_CLK_negedge or 
	 Tviol_SET_CLK_negedge or Pviol_SET or Pviol_CLK;

  VitalStateTable(
   Result => QBAR_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_ipd, QBAR_temp, D_delayed, '0', (NOT SET_ipd), CLK_delayed));
   QBAR_zd := Violation XOR  (NOT QBAR_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QBAR, true),
	             1=> (SET_ipd'last_event, tpd_SET_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFLSI_VITAL of DFFLSI is
   for VITAL_ACT
   end for;
end CFG_DFFLSI_VITAL;



 ---- CELL DFFS ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFS is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_Q		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		Q		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFS :  entity is True;
 end DFFS;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFS is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (SET_ipd,SET, tipd_SET);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, SET_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS Q_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE Q_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT SET_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFFS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_SET_CLK_posedge,
	 TimingData		=> Tmkr_SET_CLK_posedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_CLK_negedge_posedge,
	 Removal		=> thold_SET_CLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  True,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFFS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((NOT SET_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFFS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         True,
	 HeaderMsg		=> InstancePath & "DFFS",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_SET_CLK_posedge or 
	 Tviol_SET_CLK_posedge or Pviol_SET or Pviol_CLK;

  VitalStateTable(
   Result => Q_zd,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, Q_zd, D_delayed, '0', (NOT SET_ipd), CLK_ipd));
   Q_zd := Violation XOR Q_zd;
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => Q,
	 GlitchData => Q_GlitchData,
	 OutSignalName => "Q",
	 OutTemp => Q_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_Q, true),
	             1=> (SET_ipd'last_event, tpd_SET_Q, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFS_VITAL of DFFS is
   for VITAL_ACT
   end for;
end CFG_DFFS_VITAL;



 ---- CELL DFFSI ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity DFFSI is
    generic(
		TimingChecksOn: Boolean := True;
		InstancePath: String := "*";
		Xon: Boolean := False;
		MsgOn: Boolean := True;
		tpd_SET_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_CLK_QBAR		:  VitalDelayType01 := (0.100 ns, 0.100 ns);
		tsetup_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_posedge_posedge		:   VitalDelayType := 0.000 ns;
		tsetup_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_D_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		thold_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		trecovery_SET_CLK_negedge_posedge		:   VitalDelayType := 0.000 ns;
		tpw_CLK_posedge :  VitalDelayType := 0.000 ns;
		tpw_CLK_negedge  :  VitalDelayType := 0.000 ns;
		tpw_SET_posedge		:  VitalDelayType := 0.000 ns;
		tipd_SET		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_D		:   VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_CLK		:    VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		SET		:   in    STD_ULOGIC;
		CLK		:   in    STD_ULOGIC;
		D		:  in    STD_ULOGIC;
		QBAR		:  out    STD_ULOGIC);

 attribute VITAL_LEVEL0 of DFFSI :  entity is True;
 end DFFSI;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of DFFSI is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL D_ipd  : STD_ULOGIC := 'X';
	SIGNAL SET_ipd  : STD_ULOGIC := 'X';
	SIGNAL CLK_ipd : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	  VitalWireDelay (D_ipd, D, tipd_D);
	  VitalWireDelay (SET_ipd,SET, tipd_SET);
	  VitalWireDelay (CLK_ipd,CLK, tipd_CLK);
	end block;

   --------------------
   --  BEHAVIOR SECTION
   --------------------
   VITALBehavior : process (D_ipd, SET_ipd,CLK_ipd)

	-- timing check results
	VARIABLE Tviol_D_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_D_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Tviol_SET_CLK_posedge		: STD_ULOGIC := '0';
	VARIABLE Tmkr_SET_CLK_posedge		: VitalTimingDataType := VitalTimingDataInit;
	VARIABLE Pviol_CLK	: STD_ULOGIC := '0';
	VARIABLE PInfo_CLK	: VitalPeriodDataType := VitalPeriodDataInit;
	VARIABLE Pviol_SET	: STD_ULOGIC := '0';
	VARIABLE PInfo_SET	: VitalPeriodDataType := VitalPeriodDataInit;

	-- functionality results
	VARIABLE Violation	: STD_ULOGIC := '0';
	VARIABLE PrevData_Q  : STD_LOGIC_VECTOR(0 to 6);
	VARIABLE CLK_delayed	: STD_ULOGIC := 'X';
	VARIABLE D_delayed	: STD_ULOGIC := 'X';
	VARIABLE QBAR_temp	: STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS QBAR_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE QBAR_GlitchData  : VitalGlitchDataType;

   begin

   ------------------------
   --  Timing Check Section
   ------------------------
  if(TimingChecksOn) then
	VitalSetupHoldCheck (
	 Violation		=> Tviol_D_CLK_posedge,
	 TimingData		=> Tmkr_D_CLK_posedge,
	 TestSignal		=> D_ipd,
	 TestSignalName		=> "D",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName	        => "CLK",
	 RefDelay		=> 0 ns,
	 SetupHigh		=> tsetup_D_CLK_posedge_posedge,
	 SetupLow		=> tsetup_D_CLK_negedge_posedge,
	 HoldHigh		=> thold_D_CLK_posedge_posedge,
	 HoldLow		=> thold_D_CLK_negedge_posedge,
	 CheckEnabled		=>  TO_X01(((NOT SET_ipd) ) ) /= '0', 
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "/DFFSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity    => WARNING);

	VitalRecoveryRemovalCheck  (
	 Violation		=> Tviol_SET_CLK_posedge,
	 TimingData		=> Tmkr_SET_CLK_posedge,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 RefSignal		=> CLK_ipd,
	 RefSignalName		=> "CLK",
	 RefDelay		=> 0 ns,
	 Recovery		=> trecovery_SET_CLK_negedge_posedge,
	 Removal		=> thold_SET_CLK_negedge_posedge,
	 ActiveLow		 => FALSE,
	 CheckEnabled           =>  True,
	 RefTransition		=> 'R',
	 HeaderMsg		=> InstancePath & "DFFSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity	=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_CLK,
	 PeriodData		=> PInfo_CLK,
	 TestSignal		=> CLK_ipd,
	 TestSignalName		=> "CLK",
	 TestDelay		=> 0 ns,
	 Period 		=> 0 ns,
	 PulseWidthHigh		=> tpw_CLK_posedge,
	 CheckEnabled		=>		TO_X01(((NOT SET_ipd) ) ) /= '0',
	 HeaderMsg		=> InstancePath & "DFFSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	VitalPeriodPulseCheck (
	 Violation		=> Pviol_SET,
	 PeriodData		=> PInfo_SET,
	 TestSignal		=> SET_ipd,
	 TestSignalName		=> "SET",
	 TestDelay		=> 0 ns,
	 Period		=> 0 ns,
	 PulseWidthHigh		=> tpw_SET_posedge,
	 PulseWidthLow		=> 0 ns,
	 CheckEnabled		=> 			         True,
	 HeaderMsg		=> InstancePath & "DFFSI",
	 Xon		=> Xon,
	 MsgOn		=> MsgOn,
	 MsgSeverity		=> WARNING);

	end if;

	-------------------------
	--  Functionality Section
	-------------------------

	Violation := Tviol_D_CLK_posedge or 
	 Tviol_SET_CLK_posedge or 
	 Tviol_SET_CLK_posedge or Pviol_SET or Pviol_CLK;

  VitalStateTable(
   Result => QBAR_temp,
   PreviousDataIn => PrevData_Q,
   StateTable => DFEG_Q_tab,
   DataIn => (
             '1', CLK_delayed, QBAR_temp, D_delayed, '0', (NOT SET_ipd), CLK_ipd));
   QBAR_zd := Violation XOR  (NOT QBAR_temp);
   D_delayed := D_ipd;
   CLK_delayed := CLK_ipd;

	----------------------
	--  Path Delay Section
	----------------------
	VitalPathDelay01 (
	 OutSignal => QBAR,
	 GlitchData => QBAR_GlitchData,
	 OutSignalName => "QBAR",
	 OutTemp => QBAR_zd,
	 Paths => (0 => (CLK_ipd'last_event, tpd_CLK_QBAR, true),
	             1=> (SET_ipd'last_event, tpd_SET_QBAR, true)),
	 Mode => OnDetect,
	 Xon => Xon,
	 MsgOn => MsgOn,
	 MsgSeverity => WARNING);


 end process;

end VITAL_ACT;

configuration CFG_DFFSI_VITAL of DFFSI is
   for VITAL_ACT
   end for;
end CFG_DFFSI_VITAL;



 ---- CELL GLIB25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLIB25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLIB25 :  entity is True;
 end GLIB25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLIB25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);
        GL_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLIB25_VITAL of GLIB25 is 
    for VITAL_ACT
    end for;
 end CFG_GLIB25_VITAL;



 ---- CELL GLIB25LP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLIB25LP is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLIB25LP :  entity is True;
 end GLIB25LP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLIB25LP is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);
        GL_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLIB25LP_VITAL of GLIB25LP is 
    for VITAL_ACT
    end for;
 end CFG_GLIB25LP_VITAL;



 ---- CELL GLIB25LPU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLIB25LPU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLIB25LPU :  entity is True;
 end GLIB25LPU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLIB25LPU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, A_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);
        GL_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLIB25LPU_VITAL of GLIB25LPU is 
    for VITAL_ACT
    end for;
 end CFG_GLIB25LPU_VITAL;



 ---- CELL GLIB25U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLIB25U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLIB25U :  entity is True;
 end GLIB25U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLIB25U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, A_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);
        GL_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLIB25U_VITAL of GLIB25U is 
    for VITAL_ACT
    end for;
 end CFG_GLIB25U_VITAL;



 ---- CELL GLIB33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLIB33 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLIB33 :  entity is True;
 end GLIB33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLIB33 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);
        GL_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLIB33_VITAL of GLIB33 is 
    for VITAL_ACT
    end for;
 end CFG_GLIB33_VITAL;



 ---- CELL GLIB33U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLIB33U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLIB33U :  entity is True;
 end GLIB33U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLIB33U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, A_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);
        GL_zd :=TO_X01(A_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLIB33U_VITAL of GLIB33U is 
    for VITAL_ACT
    end for;
 end CFG_GLIB33U_VITAL;



 ---- CELL GLMIB25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLMIB25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLMIB25 :  entity is True;
 end GLMIB25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLMIB25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, EN_ipd, A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);
       GL_zd :=  VitalMUX2( PAD_ipd , A_ipd , (NOT EN_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true),
	             1 => (EN_ipd'last_event,tpd_EN_GL, true),
	             2 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLMIB25_VITAL of GLMIB25 is 
    for VITAL_ACT
    end for;
 end CFG_GLMIB25_VITAL;



 ---- CELL GLMIB33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLMIB33 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLMIB33 :  entity is True;
 end GLMIB33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLMIB33 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, EN_ipd, A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);
       GL_zd :=  VitalMUX2( PAD_ipd , A_ipd , (NOT EN_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true),
	             1 => (EN_ipd'last_event,tpd_EN_GL, true),
	             2 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLMIB33_VITAL of GLMIB33 is 
    for VITAL_ACT
    end for;
 end CFG_GLMIB33_VITAL;



 ---- CELL GLMIB25LP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLMIB25LP is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLMIB25LP :  entity is True;
 end GLMIB25LP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLMIB25LP is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, EN_ipd, A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);
       GL_zd :=  VitalMUX2( PAD_ipd , A_ipd , (NOT EN_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true),
	             1 => (EN_ipd'last_event,tpd_EN_GL, true),
	             2 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLMIB25LP_VITAL of GLMIB25LP is 
    for VITAL_ACT
    end for;
 end CFG_GLMIB25LP_VITAL;



 ---- CELL GLMIB25U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLMIB25U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLMIB25U :  entity is True;
 end GLMIB25U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLMIB25U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, EN_ipd, A_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);
       GL_zd :=  VitalMUX2( PAD_ipd , A_ipd , (NOT EN_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true),
	             1 => (EN_ipd'last_event,tpd_EN_GL, true),
	             2 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLMIB25U_VITAL of GLMIB25U is 
    for VITAL_ACT
    end for;
 end CFG_GLMIB25U_VITAL;



 ---- CELL GLMIB33U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLMIB33U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLMIB33U :  entity is True;
 end GLMIB33U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLMIB33U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, EN_ipd, A_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);
       GL_zd :=  VitalMUX2( PAD_ipd , A_ipd , (NOT EN_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true),
	             1 => (EN_ipd'last_event,tpd_EN_GL, true),
	             2 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLMIB33U_VITAL of GLMIB33U is 
    for VITAL_ACT
    end for;
 end CFG_GLMIB33U_VITAL;



 ---- CELL GLMIB25LPU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLMIB25LPU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLMIB25LPU :  entity is True;
 end GLMIB25LPU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLMIB25LPU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, EN_ipd, A_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);
       GL_zd :=  VitalMUX2( PAD_ipd , A_ipd , (NOT EN_ipd) );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true),
	             1 => (EN_ipd'last_event,tpd_EN_GL, true),
	             2 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLMIB25LPU_VITAL of GLMIB25LPU is 
    for VITAL_ACT
    end for;
 end CFG_GLMIB25LPU_VITAL;



 ---- CELL GLMIBL25 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLMIBL25 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLMIBL25 :  entity is True;
 end GLMIBL25;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLMIBL25 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, EN_ipd, A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);
       GL_zd :=  VitalMUX2( PAD_ipd , A_ipd , EN_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true),
	             1 => (EN_ipd'last_event,tpd_EN_GL, true),
	             2 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLMIBL25_VITAL of GLMIBL25 is 
    for VITAL_ACT
    end for;
 end CFG_GLMIBL25_VITAL;



 ---- CELL GLMIBL33 ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLMIBL33 is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLMIBL33 :  entity is True;
 end GLMIBL33;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLMIBL33 is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, EN_ipd, A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);
       GL_zd :=  VitalMUX2( PAD_ipd , A_ipd , EN_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true),
	             1 => (EN_ipd'last_event,tpd_EN_GL, true),
	             2 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLMIBL33_VITAL of GLMIBL33 is 
    for VITAL_ACT
    end for;
 end CFG_GLMIBL33_VITAL;



 ---- CELL GLMIBL25LP ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLMIBL25LP is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLMIBL25LP :  entity is True;
 end GLMIBL25LP;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLMIBL25LP is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, EN_ipd, A_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        Y_zd :=TO_X01(PAD_ipd);
       GL_zd :=  VitalMUX2( PAD_ipd , A_ipd , EN_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true),
	             1 => (EN_ipd'last_event,tpd_EN_GL, true),
	             2 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLMIBL25LP_VITAL of GLMIBL25LP is 
    for VITAL_ACT
    end for;
 end CFG_GLMIBL25LP_VITAL;



 ---- CELL GLMIBL25LPU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLMIBL25LPU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLMIBL25LPU :  entity is True;
 end GLMIBL25LPU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLMIBL25LPU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, EN_ipd, A_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);
       GL_zd :=  VitalMUX2( PAD_ipd , A_ipd , EN_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true),
	             1 => (EN_ipd'last_event,tpd_EN_GL, true),
	             2 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLMIBL25LPU_VITAL of GLMIBL25LPU is 
    for VITAL_ACT
    end for;
 end CFG_GLMIBL25LPU_VITAL;



 ---- CELL GLMIBL33U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLMIBL33U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLMIBL33U :  entity is True;
 end GLMIBL33U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLMIBL33U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, EN_ipd, A_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);
       GL_zd :=  VitalMUX2( PAD_ipd , A_ipd , EN_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true),
	             1 => (EN_ipd'last_event,tpd_EN_GL, true),
	             2 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLMIBL33U_VITAL of GLMIBL33U is 
    for VITAL_ACT
    end for;
 end CFG_GLMIBL33U_VITAL;



 ---- CELL GLMIBL25U ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity GLMIBL25U is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_PAD_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_GL		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_PAD		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		PAD		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		A		: in    STD_ULOGIC;
		Y		: out    STD_ULOGIC;
		GL		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of GLMIBL25U :  entity is True;
 end GLMIBL25U;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of GLMIBL25U is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL A_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (A_ipd, A, tipd_A);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (PAD_ipd, EN_ipd, A_ipd)


	-- functionality results
	VARIABLE PAD_ipd2 : STD_ULOGIC := 'X';
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS Y_zd : STD_LOGIC is Results(1);
	ALIAS GL_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE Y_GlitchData  : VitalGlitchDataType;
	VARIABLE GL_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
        PAD_ipd2 := VitalIdent (data => PAD_ipd,
                              ResultMap => ('U','X','0','1','H'));
        Y_zd := TO_X01(PAD_ipd2);
       GL_zd :=  VitalMUX2( PAD_ipd , A_ipd , EN_ipd );


	   ----------------------
	   --  Path Delay Section
	   ----------------------

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

     VitalPathDelay01 (
	   OutSignal => GL,
	   GlitchData => GL_GlitchData,
	   OutSignalName => "GL",
	   OutTemp => GL_zd,
	   Paths => (
	             0 => (PAD_ipd'last_event,tpd_PAD_GL, true),
	             1 => (EN_ipd'last_event,tpd_EN_GL, true),
	             2 => (A_ipd'last_event,tpd_A_GL, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_GLMIBL25U_VITAL of GLMIBL25U is 
    for VITAL_ACT
    end for;
 end CFG_GLMIBL25U_VITAL;



 ---- CELL IOB25HH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25HH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25HH :  entity is True;
 end IOB25HH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25HH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25HH_VITAL of IOB25HH is 
    for VITAL_ACT
    end for;
 end CFG_IOB25HH_VITAL;



 ---- CELL IOB25HL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25HL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25HL :  entity is True;
 end IOB25HL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25HL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25HL_VITAL of IOB25HL is 
    for VITAL_ACT
    end for;
 end CFG_IOB25HL_VITAL;



 ---- CELL IOB25HN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25HN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25HN :  entity is True;
 end IOB25HN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25HN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25HN_VITAL of IOB25HN is 
    for VITAL_ACT
    end for;
 end CFG_IOB25HN_VITAL;



 ---- CELL IOB25LH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LH :  entity is True;
 end IOB25LH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LH_VITAL of IOB25LH is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LH_VITAL;



 ---- CELL IOB25LL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LL :  entity is True;
 end IOB25LL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LL_VITAL of IOB25LL is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LL_VITAL;



 ---- CELL IOB25LN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LN :  entity is True;
 end IOB25LN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LN_VITAL of IOB25LN is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LN_VITAL;



 ---- CELL IOB25HHU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25HHU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25HHU :  entity is True;
 end IOB25HHU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25HHU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25HHU_VITAL of IOB25HHU is 
    for VITAL_ACT
    end for;
 end CFG_IOB25HHU_VITAL;



 ---- CELL IOB25HLU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25HLU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25HLU :  entity is True;
 end IOB25HLU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25HLU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25HLU_VITAL of IOB25HLU is 
    for VITAL_ACT
    end for;
 end CFG_IOB25HLU_VITAL;



 ---- CELL IOB25HNU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25HNU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25HNU :  entity is True;
 end IOB25HNU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25HNU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25HNU_VITAL of IOB25HNU is 
    for VITAL_ACT
    end for;
 end CFG_IOB25HNU_VITAL;



 ---- CELL IOB25LHU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LHU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LHU :  entity is True;
 end IOB25LHU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LHU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LHU_VITAL of IOB25LHU is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LHU_VITAL;



 ---- CELL IOB25LLU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LLU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LLU :  entity is True;
 end IOB25LLU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LLU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LLU_VITAL of IOB25LLU is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LLU_VITAL;



 ---- CELL IOB25LNU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LNU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LNU :  entity is True;
 end IOB25LNU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LNU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LNU_VITAL of IOB25LNU is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LNU_VITAL;



 ---- CELL IOB25LPHH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LPHH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LPHH :  entity is True;
 end IOB25LPHH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LPHH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LPHH_VITAL of IOB25LPHH is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LPHH_VITAL;



 ---- CELL IOB25LPHL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LPHL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LPHL :  entity is True;
 end IOB25LPHL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LPHL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LPHL_VITAL of IOB25LPHL is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LPHL_VITAL;



 ---- CELL IOB25LPHN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LPHN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LPHN :  entity is True;
 end IOB25LPHN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LPHN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LPHN_VITAL of IOB25LPHN is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LPHN_VITAL;



 ---- CELL IOB25LPLH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LPLH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LPLH :  entity is True;
 end IOB25LPLH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LPLH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LPLH_VITAL of IOB25LPLH is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LPLH_VITAL;



 ---- CELL IOB25LPLL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LPLL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LPLL :  entity is True;
 end IOB25LPLL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LPLL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LPLL_VITAL of IOB25LPLL is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LPLL_VITAL;



 ---- CELL IOB25LPLN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LPLN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LPLN :  entity is True;
 end IOB25LPLN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LPLN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LPLN_VITAL of IOB25LPLN is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LPLN_VITAL;



 ---- CELL IOB25LPHHU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LPHHU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
                tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LPHHU :  entity is True;
 end IOB25LPHHU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LPHHU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LPHHU_VITAL of IOB25LPHHU is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LPHHU_VITAL;



 ---- CELL IOB25LPHLU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LPHLU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LPHLU :  entity is True;
 end IOB25LPHLU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LPHLU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LPHLU_VITAL of IOB25LPHLU is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LPHLU_VITAL;



 ---- CELL IOB25LPHNU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LPHNU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LPHNU :  entity is True;
 end IOB25LPHNU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LPHNU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LPHNU_VITAL of IOB25LPHNU is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LPHNU_VITAL;



 ---- CELL IOB25LPLHU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LPLHU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LPLHU :  entity is True;
 end IOB25LPLHU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LPLHU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LPLHU_VITAL of IOB25LPLHU is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LPLHU_VITAL;



 ---- CELL IOB25LPLLU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LPLLU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LPLLU :  entity is True;
 end IOB25LPLLU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LPLLU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LPLLU_VITAL of IOB25LPLLU is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LPLLU_VITAL;



 ---- CELL IOB25LPLNU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB25LPLNU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB25LPLNU :  entity is True;
 end IOB25LPLNU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB25LPLNU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB25LPLNU_VITAL of IOB25LPLNU is 
    for VITAL_ACT
    end for;
 end CFG_IOB25LPLNU_VITAL;



 ---- CELL IOB33LH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB33LH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB33LH :  entity is True;
 end IOB33LH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB33LH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB33LH_VITAL of IOB33LH is 
    for VITAL_ACT
    end for;
 end CFG_IOB33LH_VITAL;



 ---- CELL IOB33LL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB33LL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB33LL :  entity is True;
 end IOB33LL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB33LL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB33LL_VITAL of IOB33LL is 
    for VITAL_ACT
    end for;
 end CFG_IOB33LL_VITAL;



 ---- CELL IOB33LN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB33LN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB33LN :  entity is True;
 end IOB33LN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB33LN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB33LN_VITAL of IOB33LN is 
    for VITAL_ACT
    end for;
 end CFG_IOB33LN_VITAL;



 ---- CELL IOB33PH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB33PH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB33PH :  entity is True;
 end IOB33PH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB33PH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB33PH_VITAL of IOB33PH is 
    for VITAL_ACT
    end for;
 end CFG_IOB33PH_VITAL;



 ---- CELL IOB33PL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB33PL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB33PL :  entity is True;
 end IOB33PL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB33PL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB33PL_VITAL of IOB33PL is 
    for VITAL_ACT
    end for;
 end CFG_IOB33PL_VITAL;



 ---- CELL IOB33PN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB33PN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB33PN :  entity is True;
 end IOB33PN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB33PN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB33PN_VITAL of IOB33PN is 
    for VITAL_ACT
    end for;
 end CFG_IOB33PN_VITAL;



 ---- CELL IOB33LHU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB33LHU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB33LHU :  entity is True;
 end IOB33LHU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB33LHU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB33LHU_VITAL of IOB33LHU is 
    for VITAL_ACT
    end for;
 end CFG_IOB33LHU_VITAL;



 ---- CELL IOB33LLU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB33LLU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB33LLU :  entity is True;
 end IOB33LLU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB33LLU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB33LLU_VITAL of IOB33LLU is 
    for VITAL_ACT
    end for;
 end CFG_IOB33LLU_VITAL;



 ---- CELL IOB33LNU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB33LNU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB33LNU :  entity is True;
 end IOB33LNU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB33LNU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB33LNU_VITAL of IOB33LNU is 
    for VITAL_ACT
    end for;
 end CFG_IOB33LNU_VITAL;



 ---- CELL IOB33PHU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB33PHU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB33PHU :  entity is True;
 end IOB33PHU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB33PHU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB33PHU_VITAL of IOB33PHU is 
    for VITAL_ACT
    end for;
 end CFG_IOB33PHU_VITAL;



 ---- CELL IOB33PLU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB33PLU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB33PLU :  entity is True;
 end IOB33PLU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB33PLU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB33PLU_VITAL of IOB33PLU is 
    for VITAL_ACT
    end for;
 end CFG_IOB33PLU_VITAL;



 ---- CELL IOB33PNU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOB33PNU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOB33PNU :  entity is True;
 end IOB33PNU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOB33PNU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOB33PNU_VITAL of IOB33PNU is 
    for VITAL_ACT
    end for;
 end CFG_IOB33PNU_VITAL;



 ---- CELL IOBL25HH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25HH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25HH :  entity is True;
 end IOBL25HH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25HH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25HH_VITAL of IOBL25HH is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25HH_VITAL;



 ---- CELL IOBL25HL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25HL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25HL :  entity is True;
 end IOBL25HL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25HL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25HL_VITAL of IOBL25HL is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25HL_VITAL;



 ---- CELL IOBL25HN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25HN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25HN :  entity is True;
 end IOBL25HN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25HN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25HN_VITAL of IOBL25HN is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25HN_VITAL;



 ---- CELL IOBL25LH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LH :  entity is True;
 end IOBL25LH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LH_VITAL of IOBL25LH is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LH_VITAL;



 ---- CELL IOBL25LL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LL :  entity is True;
 end IOBL25LL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LL_VITAL of IOBL25LL is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LL_VITAL;



 ---- CELL IOBL25LN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LN :  entity is True;
 end IOBL25LN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LN_VITAL of IOBL25LN is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LN_VITAL;



 ---- CELL IOBL25HHU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25HHU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25HHU :  entity is True;
 end IOBL25HHU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25HHU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25HHU_VITAL of IOBL25HHU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25HHU_VITAL;



 ---- CELL IOBL25HLU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25HLU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25HLU :  entity is True;
 end IOBL25HLU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25HLU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25HLU_VITAL of IOBL25HLU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25HLU_VITAL;



 ---- CELL IOBL25HNU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25HNU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25HNU :  entity is True;
 end IOBL25HNU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25HNU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25HNU_VITAL of IOBL25HNU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25HNU_VITAL;



 ---- CELL IOBL25LHU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LHU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LHU :  entity is True;
 end IOBL25LHU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LHU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LHU_VITAL of IOBL25LHU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LHU_VITAL;



 ---- CELL IOBL25LLU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LLU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LLU :  entity is True;
 end IOBL25LLU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LLU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LLU_VITAL of IOBL25LLU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LLU_VITAL;



 ---- CELL IOBL25LNU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LNU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LNU :  entity is True;
 end IOBL25LNU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LNU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LNU_VITAL of IOBL25LNU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LNU_VITAL;



 ---- CELL IOBL25LPHH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LPHH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LPHH :  entity is True;
 end IOBL25LPHH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LPHH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LPHH_VITAL of IOBL25LPHH is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LPHH_VITAL;



 ---- CELL IOBL25LPHL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LPHL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LPHL :  entity is True;
 end IOBL25LPHL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LPHL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LPHL_VITAL of IOBL25LPHL is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LPHL_VITAL;



 ---- CELL IOBL25LPHN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LPHN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LPHN :  entity is True;
 end IOBL25LPHN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LPHN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LPHN_VITAL of IOBL25LPHN is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LPHN_VITAL;



 ---- CELL IOBL25LPLH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LPLH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LPLH :  entity is True;
 end IOBL25LPLH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LPLH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LPLH_VITAL of IOBL25LPLH is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LPLH_VITAL;



 ---- CELL IOBL25LPLL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LPLL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LPLL :  entity is True;
 end IOBL25LPLL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LPLL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LPLL_VITAL of IOBL25LPLL is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LPLL_VITAL;



 ---- CELL IOBL25LPLN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LPLN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LPLN :  entity is True;
 end IOBL25LPLN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LPLN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LPLN_VITAL of IOBL25LPLN is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LPLN_VITAL;



 ---- CELL IOBL25LPHHU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LPHHU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LPHHU :  entity is True;
 end IOBL25LPHHU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LPHHU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LPHHU_VITAL of IOBL25LPHHU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LPHHU_VITAL;



 ---- CELL IOBL25LPHLU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LPHLU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LPHLU :  entity is True;
 end IOBL25LPHLU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LPHLU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LPHLU_VITAL of IOBL25LPHLU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LPHLU_VITAL;



 ---- CELL IOBL25LPHNU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LPHNU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LPHNU :  entity is True;
 end IOBL25LPHNU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LPHNU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LPHNU_VITAL of IOBL25LPHNU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LPHNU_VITAL;



 ---- CELL IOBL25LPLHU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LPLHU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LPLHU :  entity is True;
 end IOBL25LPLHU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LPLHU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LPLHU_VITAL of IOBL25LPLHU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LPLHU_VITAL;



 ---- CELL IOBL25LPLLU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LPLLU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LPLLU :  entity is True;
 end IOBL25LPLLU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LPLLU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LPLLU_VITAL of IOBL25LPLLU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LPLLU_VITAL;



 ---- CELL IOBL25LPLNU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL25LPLNU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL25LPLNU :  entity is True;
 end IOBL25LPLNU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL25LPLNU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL25LPLNU_VITAL of IOBL25LPLNU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL25LPLNU_VITAL;



 ---- CELL IOBL33LH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL33LH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL33LH :  entity is True;
 end IOBL33LH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL33LH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL33LH_VITAL of IOBL33LH is 
    for VITAL_ACT
    end for;
 end CFG_IOBL33LH_VITAL;



 ---- CELL IOBL33LL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL33LL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL33LL :  entity is True;
 end IOBL33LL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL33LL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL33LL_VITAL of IOBL33LL is 
    for VITAL_ACT
    end for;
 end CFG_IOBL33LL_VITAL;



 ---- CELL IOBL33LN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL33LN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL33LN :  entity is True;
 end IOBL33LN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL33LN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL33LN_VITAL of IOBL33LN is 
    for VITAL_ACT
    end for;
 end CFG_IOBL33LN_VITAL;



 ---- CELL IOBL33PH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL33PH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL33PH :  entity is True;
 end IOBL33PH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL33PH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL33PH_VITAL of IOBL33PH is 
    for VITAL_ACT
    end for;
 end CFG_IOBL33PH_VITAL;



 ---- CELL IOBL33PL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL33PL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL33PL :  entity is True;
 end IOBL33PL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL33PL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL33PL_VITAL of IOBL33PL is 
    for VITAL_ACT
    end for;
 end CFG_IOBL33PL_VITAL;



 ---- CELL IOBL33PN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL33PN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL33PN :  entity is True;
 end IOBL33PN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL33PN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL33PN_VITAL of IOBL33PN is 
    for VITAL_ACT
    end for;
 end CFG_IOBL33PN_VITAL;



 ---- CELL IOBL33LHU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL33LHU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL33LHU :  entity is True;
 end IOBL33LHU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL33LHU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL33LHU_VITAL of IOBL33LHU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL33LHU_VITAL;



 ---- CELL IOBL33LLU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL33LLU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL33LLU :  entity is True;
 end IOBL33LLU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL33LLU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL33LLU_VITAL of IOBL33LLU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL33LLU_VITAL;



 ---- CELL IOBL33LNU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL33LNU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL33LNU :  entity is True;
 end IOBL33LNU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL33LNU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL33LNU_VITAL of IOBL33LNU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL33LNU_VITAL;



 ---- CELL IOBL33PHU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL33PHU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL33PHU :  entity is True;
 end IOBL33PHU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL33PHU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL33PHU_VITAL of IOBL33PHU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL33PHU_VITAL;



 ---- CELL IOBL33PLU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL33PLU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL33PLU :  entity is True;
 end IOBL33PLU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL33PLU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL33PLU_VITAL of IOBL33PLU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL33PLU_VITAL;



 ---- CELL IOBL33PNU ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity IOBL33PNU is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tpd_PAD_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_A_Y		: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_Y	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_PAD	: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: inout STD_ULOGIC;
		Y		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of IOBL33PNU :  entity is True;
 end IOBL33PNU;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of IOBL33PNU is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';
	SIGNAL PAD_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	VitalWireDelay (PAD_ipd, PAD, tipd_PAD);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd, PAD_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 2)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);
	ALIAS Y_zd : STD_LOGIC is Results(2);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;
	VARIABLE Y_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);
        Y_zd :=TO_X01(PAD_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01HWLH-");

     VitalPathDelay01 (
	   OutSignal => Y,
	   GlitchData => Y_GlitchData,
	   OutSignalName => "Y",
	   OutTemp => Y_zd,
	   Paths => (
	             0 => (A_ipd'last_event,tpd_A_Y, true),
	             1 => (EN_ipd'last_event,tpd_EN_Y, true),
	             2 => (PAD_ipd'last_event,tpd_PAD_Y, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING);

 end process;

end VITAL_ACT;

 configuration CFG_IOBL33PNU_VITAL of IOBL33PNU is 
    for VITAL_ACT
    end for;
 end CFG_IOBL33PNU_VITAL;



 ---- CELL OTB25HH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB25HH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB25HH :  entity is True;
 end OTB25HH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB25HH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB25HH_VITAL of OTB25HH is 
    for VITAL_ACT
    end for;
 end CFG_OTB25HH_VITAL;



 ---- CELL OTB25HL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB25HL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB25HL :  entity is True;
 end OTB25HL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB25HL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB25HL_VITAL of OTB25HL is 
    for VITAL_ACT
    end for;
 end CFG_OTB25HL_VITAL;



 ---- CELL OTB25HN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB25HN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB25HN :  entity is True;
 end OTB25HN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB25HN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB25HN_VITAL of OTB25HN is 
    for VITAL_ACT
    end for;
 end CFG_OTB25HN_VITAL;



 ---- CELL OTB25LH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB25LH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB25LH :  entity is True;
 end OTB25LH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB25LH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB25LH_VITAL of OTB25LH is 
    for VITAL_ACT
    end for;
 end CFG_OTB25LH_VITAL;



 ---- CELL OTB25LL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB25LL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB25LL :  entity is True;
 end OTB25LL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB25LL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB25LL_VITAL of OTB25LL is 
    for VITAL_ACT
    end for;
 end CFG_OTB25LL_VITAL;



 ---- CELL OTB25LN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB25LN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB25LN :  entity is True;
 end OTB25LN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB25LN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB25LN_VITAL of OTB25LN is 
    for VITAL_ACT
    end for;
 end CFG_OTB25LN_VITAL;



 ---- CELL OTB25LPLH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB25LPLH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB25LPLH :  entity is True;
 end OTB25LPLH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB25LPLH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB25LPLH_VITAL of OTB25LPLH is 
    for VITAL_ACT
    end for;
 end CFG_OTB25LPLH_VITAL;



 ---- CELL OTB25LPLL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB25LPLL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB25LPLL :  entity is True;
 end OTB25LPLL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB25LPLL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB25LPLL_VITAL of OTB25LPLL is 
    for VITAL_ACT
    end for;
 end CFG_OTB25LPLL_VITAL;



 ---- CELL OTB25LPLN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB25LPLN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB25LPLN :  entity is True;
 end OTB25LPLN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB25LPLN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB25LPLN_VITAL of OTB25LPLN is 
    for VITAL_ACT
    end for;
 end CFG_OTB25LPLN_VITAL;



 ---- CELL OTB25LPHH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB25LPHH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB25LPHH :  entity is True;
 end OTB25LPHH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB25LPHH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB25LPHH_VITAL of OTB25LPHH is 
    for VITAL_ACT
    end for;
 end CFG_OTB25LPHH_VITAL;



 ---- CELL OTB25LPHL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB25LPHL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB25LPHL :  entity is True;
 end OTB25LPHL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB25LPHL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB25LPHL_VITAL of OTB25LPHL is 
    for VITAL_ACT
    end for;
 end CFG_OTB25LPHL_VITAL;



 ---- CELL OTB25LPHN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB25LPHN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB25LPHN :  entity is True;
 end OTB25LPHN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB25LPHN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB25LPHN_VITAL of OTB25LPHN is 
    for VITAL_ACT
    end for;
 end CFG_OTB25LPHN_VITAL;



 ---- CELL OTB33LH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB33LH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB33LH :  entity is True;
 end OTB33LH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB33LH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB33LH_VITAL of OTB33LH is 
    for VITAL_ACT
    end for;
 end CFG_OTB33LH_VITAL;



 ---- CELL OTB33LL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB33LL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB33LL :  entity is True;
 end OTB33LL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB33LL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB33LL_VITAL of OTB33LL is 
    for VITAL_ACT
    end for;
 end CFG_OTB33LL_VITAL;



 ---- CELL OTB33LN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB33LN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB33LN :  entity is True;
 end OTB33LN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB33LN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB33LN_VITAL of OTB33LN is 
    for VITAL_ACT
    end for;
 end CFG_OTB33LN_VITAL;



 ---- CELL OTB33PH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB33PH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB33PH :  entity is True;
 end OTB33PH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB33PH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB33PH_VITAL of OTB33PH is 
    for VITAL_ACT
    end for;
 end CFG_OTB33PH_VITAL;



 ---- CELL OTB33PL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB33PL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB33PL :  entity is True;
 end OTB33PL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB33PL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB33PL_VITAL of OTB33PL is 
    for VITAL_ACT
    end for;
 end CFG_OTB33PL_VITAL;



 ---- CELL OTB33PN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTB33PN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTB33PN :  entity is True;
 end OTB33PN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTB33PN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>(NOT EN_ipd));


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTB33PN_VITAL of OTB33PN is 
    for VITAL_ACT
    end for;
 end CFG_OTB33PN_VITAL;



 ---- CELL OTBL25HH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL25HH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL25HH :  entity is True;
 end OTBL25HH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL25HH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL25HH_VITAL of OTBL25HH is 
    for VITAL_ACT
    end for;
 end CFG_OTBL25HH_VITAL;



 ---- CELL OTBL25HL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL25HL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL25HL :  entity is True;
 end OTBL25HL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL25HL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL25HL_VITAL of OTBL25HL is 
    for VITAL_ACT
    end for;
 end CFG_OTBL25HL_VITAL;



 ---- CELL OTBL25HN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL25HN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL25HN :  entity is True;
 end OTBL25HN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL25HN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL25HN_VITAL of OTBL25HN is 
    for VITAL_ACT
    end for;
 end CFG_OTBL25HN_VITAL;



 ---- CELL OTBL25LH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL25LH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL25LH :  entity is True;
 end OTBL25LH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL25LH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL25LH_VITAL of OTBL25LH is 
    for VITAL_ACT
    end for;
 end CFG_OTBL25LH_VITAL;



 ---- CELL OTBL25LL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL25LL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL25LL :  entity is True;
 end OTBL25LL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL25LL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL25LL_VITAL of OTBL25LL is 
    for VITAL_ACT
    end for;
 end CFG_OTBL25LL_VITAL;



 ---- CELL OTBL25LN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL25LN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL25LN :  entity is True;
 end OTBL25LN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL25LN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL25LN_VITAL of OTBL25LN is 
    for VITAL_ACT
    end for;
 end CFG_OTBL25LN_VITAL;



 ---- CELL OTBL25LPLH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL25LPLH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL25LPLH :  entity is True;
 end OTBL25LPLH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL25LPLH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL25LPLH_VITAL of OTBL25LPLH is 
    for VITAL_ACT
    end for;
 end CFG_OTBL25LPLH_VITAL;



 ---- CELL OTBL25LPLL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL25LPLL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL25LPLL :  entity is True;
 end OTBL25LPLL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL25LPLL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL25LPLL_VITAL of OTBL25LPLL is 
    for VITAL_ACT
    end for;
 end CFG_OTBL25LPLL_VITAL;



 ---- CELL OTBL25LPLN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL25LPLN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL25LPLN :  entity is True;
 end OTBL25LPLN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL25LPLN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL25LPLN_VITAL of OTBL25LPLN is 
    for VITAL_ACT
    end for;
 end CFG_OTBL25LPLN_VITAL;



 ---- CELL OTBL25LPHH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL25LPHH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL25LPHH :  entity is True;
 end OTBL25LPHH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL25LPHH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL25LPHH_VITAL of OTBL25LPHH is 
    for VITAL_ACT
    end for;
 end CFG_OTBL25LPHH_VITAL;



 ---- CELL OTBL25LPHL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL25LPHL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL25LPHL :  entity is True;
 end OTBL25LPHL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL25LPHL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL25LPHL_VITAL of OTBL25LPHL is 
    for VITAL_ACT
    end for;
 end CFG_OTBL25LPHL_VITAL;



 ---- CELL OTBL25LPHN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL25LPHN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL25LPHN :  entity is True;
 end OTBL25LPHN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL25LPHN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL25LPHN_VITAL of OTBL25LPHN is 
    for VITAL_ACT
    end for;
 end CFG_OTBL25LPHN_VITAL;



 ---- CELL OTBL33LH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL33LH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL33LH :  entity is True;
 end OTBL33LH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL33LH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL33LH_VITAL of OTBL33LH is 
    for VITAL_ACT
    end for;
 end CFG_OTBL33LH_VITAL;



 ---- CELL OTBL33LL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL33LL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL33LL :  entity is True;
 end OTBL33LL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL33LL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL33LL_VITAL of OTBL33LL is 
    for VITAL_ACT
    end for;
 end CFG_OTBL33LL_VITAL;



 ---- CELL OTBL33LN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL33LN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL33LN :  entity is True;
 end OTBL33LN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL33LN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL33LN_VITAL of OTBL33LN is 
    for VITAL_ACT
    end for;
 end CFG_OTBL33LN_VITAL;



 ---- CELL OTBL33PH ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL33PH is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL33PH :  entity is True;
 end OTBL33PH;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL33PH is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL33PH_VITAL of OTBL33PH is 
    for VITAL_ACT
    end for;
 end CFG_OTBL33PH_VITAL;



 ---- CELL OTBL33PL ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL33PL is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL33PL :  entity is True;
 end OTBL33PL;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL33PL is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL33PL_VITAL of OTBL33PL is 
    for VITAL_ACT
    end for;
 end CFG_OTBL33PL_VITAL;



 ---- CELL OTBL33PN ----
 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 library IEEE;
 use IEEE.VITAL_Timing.all;

 ---- entity declaration ----
 entity OTBL33PN is
    generic(
		TimingChecksOn:Boolean := True;
		Xon: Boolean := False;
		InstancePath: String :="*";
		MsgOn: Boolean := True;
		tpd_A_PAD	: VitalDelayType01 := (0.100 ns, 0.100 ns);
		tpd_EN_PAD : VitalDelayType01z := (0.0 ns, 0.0 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
		tipd_A		: VitalDelayType01 := (0.000 ns, 0.000 ns);
		tipd_EN		: VitalDelayType01 := (0.000 ns, 0.000 ns));


    port(
		A		: in    STD_ULOGIC;
		EN		: in    STD_ULOGIC;
		PAD		: out    STD_ULOGIC);
 attribute VITAL_LEVEL0 of OTBL33PN :  entity is True;
 end OTBL33PN;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
library a500k;
use a500k.VTABLES.all;

architecture VITAL_ACT of OTBL33PN is
	attribute VITAL_LEVEL1 of VITAL_ACT : architecture is True;

	SIGNAL A_ipd  : STD_ULOGIC := 'X';
	SIGNAL EN_ipd  : STD_ULOGIC := 'X';

begin

	---------------------
	--  INPUT PATH DELAYs
	---------------------
	WireDelay : block
	begin
	VitalWireDelay (A_ipd, A, tipd_A);
	VitalWireDelay (EN_ipd, EN, tipd_EN);
	end block;

	--------------------
	--  BEHAVIOR SECTION
	--------------------
	VITALBehavior : process (A_ipd, EN_ipd)


	-- functionality results
	VARIABLE Results : STD_LOGIC_VECTOR(1 to 1)  := (others => 'X');
	ALIAS PAD_zd : STD_LOGIC is Results(1);

	-- output glitch detection variables
	VARIABLE PAD_GlitchData  : VitalGlitchDataType;

	begin

	   -------------------------
	   --  Functionality Section
	   -------------------------
       PAD_zd := VitalBUFIF0 (data => A_ipd,
                   enable =>EN_ipd);


	   ----------------------
	   --  Path Delay Section
	   ----------------------

	  VitalPathDelay01Z (
	   OutSignal => PAD,
	   GlitchData => PAD_GlitchData,
	   OutSignalName => "PAD",
	   OutTemp => PAD_zd,
	   Paths => (
	             0 => (A_ipd'last_event,VitalExtendToFillDelay(tpd_A_PAD),true),
	             1 => (EN_ipd'last_event,tpd_EN_PAD, true)),
	  Mode => OnDetect,
	  Xon => Xon,
	  MsgOn => MsgOn,
	  MsgSeverity => WARNING,
	  OutputMap => "UX01ZWLH-");

 end process;

end VITAL_ACT;

 configuration CFG_OTBL33PN_VITAL of OTBL33PN is 
    for VITAL_ACT
    end for;
 end CFG_OTBL33PN_VITAL;


----------------------------------------------------------------------- 
--   ACTEL A500K UJTAG VITAL Model
--
--   Revision 1.1 -  9/17/03.
-----------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
library IEEE;
use IEEE.VITAL_Timing.all;

-- entity declaration --
entity UJTAG is
   generic(
      TimingChecksOn : Boolean := True;
      InstancePath   : String  := "*";
      Xon            : Boolean := False;
      MsgOn          : Boolean := True;

      tipd_UTDO      : VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_TMS       : VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_TDI       : VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_TCK       : VitalDelayType01 := (0.0 ns, 0.0 ns);
      tipd_TRSTB     : VitalDelayType01 := (0.0 ns, 0.0 ns)
     );

   port(
      UTDO           :	in    STD_ULOGIC; 
      TMS            :	in    STD_ULOGIC;
      TDI            :	in    STD_ULOGIC;  
      TCK            :	in    STD_ULOGIC;
      TRSTB          :	in    STD_ULOGIC; 
      UIREG0         :  out   STD_ULOGIC;
      UIREG1         :  out   STD_ULOGIC;
      UIREG2         :  out   STD_ULOGIC;
      UIREG3         :  out   STD_ULOGIC;
      UIREG4         :  out   STD_ULOGIC;
      UIREG5         :  out   STD_ULOGIC;
      UIREG6         :  out   STD_ULOGIC;
      UIREG7         :  out   STD_ULOGIC;
      UTDI           :  out   STD_ULOGIC;
      URSTB          :  out   STD_ULOGIC;
      UDRCK          :  out   STD_ULOGIC;
      UDRSH          :  out   STD_ULOGIC;
      UDRUPD         :  out   STD_ULOGIC;
      TDO            :  out   STD_ULOGIC);            

  attribute VITAL_LEVEL0 of UJTAG : entity is True;
end UJTAG;

-- architecture body --
library IEEE;
use IEEE.VITAL_Primitives.all;
architecture VITAL_ACT of UJTAG is
   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   SIGNAL UTDO_ipd          : STD_ULOGIC := 'X';
   SIGNAL TMS_ipd           : STD_ULOGIC := 'X';
   SIGNAL TDI_ipd           : STD_ULOGIC := 'X';
   SIGNAL TCK_ipd           : STD_ULOGIC := 'X';
   SIGNAL TRSTB_ipd         : STD_ULOGIC := 'X';

   SIGNAL SHREG             : std_logic_vector(7 downto 0) := "XXXXXXXX";
   SIGNAL IR                : std_logic_vector(7 downto 0);

   type state_type is (Test_Logic_Reset,
                       Run_Test_Idle,
                       Select_DR,
                       Capture_DR,
                       Shift_DR,
                       Exit1_DR,
                       Pause_DR,
                       Exit2_DR,
                       Update_DR,
                       Select_IR,
                       Capture_IR,
                       Shift_IR,
                       Exit1_IR,
                       Pause_IR,
                       Exit2_IR,
                       Update_IR,
                       Unknown
                      );

   SIGNAL STATE : state_type := Unknown;

begin

   ---------------------
   --  INPUT PATH DELAYs
   ---------------------
   WireDelay : block

   begin

     VitalWireDelay (UTDO_ipd, UTDO, tipd_UTDO);
     VitalWireDelay (TMS_ipd, TMS, tipd_TMS);
     VitalWireDelay (TDI_ipd, TDI, tipd_TDI);
     VitalWireDelay (TCK_ipd, TCK, tipd_TCK);
     VitalWireDelay (TRSTB_ipd, TRSTB, tipd_TRSTB);

   end block WireDelay;

  -- #########################################################
  -- # Behavior Section
  -- #########################################################

  OUTPUTS1 : process (TCK_ipd, TRSTB_ipd)

  begin
    if ((TRSTB_ipd'event) and (TO_X01(TRSTB_ipd) = '0')) then
                UDRUPD <= '0';
                UDRSH  <= '0';
  
    elsif ((TCK_ipd'event) and (TO_X01(TCK_ipd) = '0')) then
      if (STATE = Unknown) then
        UDRUPD <= 'X';
        UDRSH  <= 'X';
      else
        if (STATE = Update_DR) then
          UDRUPD <= '1';
        else
          UDRUPD <= '0';
        end if;
    
        if (STATE = Shift_DR) then
          UDRSH  <= '1';
        else
          UDRSH  <= '0';
        end if;

      end if;
    end if;

  end process OUTPUTS1;

  STATES: process (TCK_ipd, TRSTB_ipd)
  begin
    if ((TRSTB_ipd'event) and (TO_X01(TRSTB_ipd) = '0')) then
       STATE <= Test_Logic_Reset;
    elsif ((TCK_ipd'event) and (TO_X01(TCK_ipd) = '1')) then
       case STATE is
         when Test_Logic_Reset       => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Test_Logic_Reset;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Run_Test_Idle;
                                        end if;
         when Run_Test_Idle          => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Select_DR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Run_Test_Idle;
                                        end if;
         when Select_DR              => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Select_IR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Capture_DR;
                                        end if;
         when Capture_DR | Shift_DR  => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Exit1_DR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Shift_DR;
                                        end if;
         when Exit1_DR               => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Update_DR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Pause_DR;
                                        end if;
         when Pause_DR               => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Exit2_DR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Pause_DR;
                                        end if;
         when Exit2_DR               => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Update_DR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Shift_DR;
                                        end if;
         when  Select_IR             => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Test_Logic_Reset;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Capture_IR;
                                        end if;
         when Capture_IR | Shift_IR  => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Exit1_IR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Shift_IR;
                                        end if;
         when Exit1_IR               => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Update_IR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Pause_IR;
                                        end if;
         when Pause_IR               => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <=  Exit2_IR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Pause_IR;
                                        end if;
         when Exit2_IR               => if (TO_X01(TMS_ipd) = '1') then
                                          STATE <= Update_IR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Shift_IR;
                                        end if;
         when Update_DR | Update_IR  => if (TO_X01(TMS_ipd)= '1') then
                                          STATE <= Select_DR;
                                        elsif (TO_X01(TMS_ipd) = '0') then
                                          STATE <= Run_Test_Idle;
                                        end if;
         when Unknown                => STATE <= Unknown;
       end case;
    end if;
  end process STATES;

  CLOCK_SHREG: process(TCK_ipd)
  begin
    if ((TCK_ipd'event) and (TO_X01(TCK_ipd) = '1')) then
      case STATE is
        when Capture_IR  => SHREG <=  "XXXXXX01";
        when Capture_DR  => SHREG <=  "00000000";
        when Shift_IR | Shift_DR  => SHREG <= TDI_ipd & SHREG(7) & SHREG(6) & SHREG(5) 
                                              & SHREG(4) & SHREG(3) & SHREG(2) & SHREG(1);
    
        when others   => SHREG <= SHREG;  
      end case;
    end if;
  end process CLOCK_SHREG;


  OUTPUTS2: process(TCK_ipd, TRSTB_ipd)
  begin
    if ((TRSTB_ipd'event) and (TO_X01(TRSTB_ipd) = '0')) then
      IR <= "11111111"; -- Bypass
      TDO <= 'Z';
    elsif ((TCK_ipd'event) and (TO_X01(TCK_ipd) = '0')) then
      if (STATE = Shift_IR) then
        TDO <= SHREG(0);
      elsif (STATE = Shift_DR) then
        if (IR(7) = '0' and (IR(6) = '1' or IR(5) = '1' or IR(4) = '1')) then
          TDO <= UTDO;
        else
          TDO <= SHREG(7);
        end if;
      elsif (STATE = Update_IR) then
        TDO <= 'Z';
        IR <= SHREG;
      else
        TDO <= 'Z';
      end if;
    end if;
  end process OUTPUTS2;

  OUTPUTS3: process(IR)
  begin
    UIREG7 <= IR(7);
    UIREG6 <= IR(6);
    UIREG5 <= IR(5);
    UIREG4 <= IR(4);
    UIREG3 <= IR(3);
    UIREG2 <= IR(2);
    UIREG1 <= IR(1);
    UIREG0 <= IR(0);
  end process OUTPUTS3;

--  OUTPUTS4: process(TDI_ipd)
--  begin
--    UTDI <= TDI_ipd;
--  end process;

UTDI <= TDI_ipd;

  OUTPUTS5: process(TCK_ipd, STATE)
  begin
    if (TO_X01(TCK_ipd) = 'X') then 
      UDRCK <= 'X';
    elsif (TO_X01(TCK_ipd) = '1') then 
      UDRCK <= '1';
    elsif (STATE = Unknown) then
      UDRCK <= 'X';
    elsif (STATE /= Shift_DR and STATE /= Capture_DR) then
      UDRCK <= '1';
    else
      UDRCK <= '0';
    end if;
  end process;

  OUTPUTS6: process(STATE)
  begin
    if (STATE = Unknown) then
      URSTB <= 'X';
    elsif (STATE = Test_Logic_Reset) then
      URSTB <= '0';
    else
      URSTB <= '1';
    end if;
  end process;

       
end VITAL_ACT;

configuration CFG_UJTAG_VITAL of UJTAG is
  for VITAL_ACT
  end for;
end CFG_UJTAG_VITAL;


---- CELL RAM256x9AA ----

LIBRARY ieee;
LIBRARY STD;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

USE std.textio.all;
USE ieee.std_logic_textio.all;
LIBRARY a500k;
USE a500k.all;

entity RAM256x9AA is 

   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI0_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI1_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI2_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI3_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI4_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI5_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI6_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI7_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI8_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns,0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpw_RDB_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_RDB_negedge	        : VitalDelayType := 0.000 ns;
 	tperiod_RDB	        : VitalDelayType := 0.000 ns;
 	tpw_RBLKB_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RBLKB_negedge	: VitalDelayType := 0.000 ns;
 	tperiod_RBLKB	        : VitalDelayType := 0.000 ns;
 	tpw_RADDR0_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR0_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                           : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                         : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                         : VitalDelayType := 0.000 ns;
 	tperiod_WRB                             : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_RDB_WRB_negedge_negedge          : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_WRB_posedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RBLKB_WRB_posedge_posedge         : VitalDelayType := 0.000 ns;
 	thold_RDB_WBLKB_posedge_posedge         : VitalDelayType := 0.000 ns;
 	thold_RBLKB_WBLKB_posedge_posedge       : VitalDelayType := 0.000 ns;
 	thold_RADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';
   WPE    :  OUT STD_LOGIC := 'X';
   RPE    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');

ATTRIBUTE VITAL_LEVEL0 OF RAM256x9AA : entity IS True ;
END RAM256x9AA;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of RAM256x9AA is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal WADDR0_ipd : std_ulogic := 'X';
   signal WADDR1_ipd : std_ulogic := 'X';
   signal WADDR2_ipd : std_ulogic := 'X';
   signal WADDR3_ipd : std_ulogic := 'X';
   signal WADDR4_ipd : std_ulogic := 'X';
   signal WADDR5_ipd : std_ulogic := 'X';
   signal WADDR6_ipd : std_ulogic := 'X';
   signal WADDR7_ipd : std_ulogic := 'X';
   signal RADDR0_ipd : std_ulogic := 'X';
   signal RADDR1_ipd : std_ulogic := 'X';
   signal RADDR2_ipd : std_ulogic := 'X';
   signal RADDR3_ipd : std_ulogic := 'X';
   signal RADDR4_ipd : std_ulogic := 'X';
   signal RADDR5_ipd : std_ulogic := 'X';
   signal RADDR6_ipd : std_ulogic := 'X';
   signal RADDR7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

	-- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';
   signal INIT_MEM   : std_logic:= '0';
   signal WBdlyd     : std_ulogic := 'X';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic:= 'X';
   signal par_f2     : std_logic:= 'X';

 begin  --  VITAL_ACT
   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (WADDR0_ipd, WADDR0, VitalExtendToFillDelay(tipd_WADDR0));
   VitalWireDelay (WADDR1_ipd, WADDR1, VitalExtendToFillDelay(tipd_WADDR1));
   VitalWireDelay (WADDR2_ipd, WADDR2, VitalExtendToFillDelay(tipd_WADDR2));
   VitalWireDelay (WADDR3_ipd, WADDR3, VitalExtendToFillDelay(tipd_WADDR3));
   VitalWireDelay (WADDR4_ipd, WADDR4, VitalExtendToFillDelay(tipd_WADDR4));
   VitalWireDelay (WADDR5_ipd, WADDR5, VitalExtendToFillDelay(tipd_WADDR5));
   VitalWireDelay (WADDR6_ipd, WADDR6, VitalExtendToFillDelay(tipd_WADDR6));
   VitalWireDelay (WADDR7_ipd, WADDR7, VitalExtendToFillDelay(tipd_WADDR7));
   VitalWireDelay (RADDR0_ipd, RADDR0, VitalExtendToFillDelay(tipd_RADDR0));
   VitalWireDelay (RADDR1_ipd, RADDR1, VitalExtendToFillDelay(tipd_RADDR1));
   VitalWireDelay (RADDR2_ipd, RADDR2, VitalExtendToFillDelay(tipd_RADDR2));
   VitalWireDelay (RADDR3_ipd, RADDR3, VitalExtendToFillDelay(tipd_RADDR3));
   VitalWireDelay (RADDR4_ipd, RADDR4, VitalExtendToFillDelay(tipd_RADDR4));
   VitalWireDelay (RADDR5_ipd, RADDR5, VitalExtendToFillDelay(tipd_RADDR5));
   VitalWireDelay (RADDR6_ipd, RADDR6, VitalExtendToFillDelay(tipd_RADDR6));
   VitalWireDelay (RADDR7_ipd, RADDR7, VitalExtendToFillDelay(tipd_RADDR7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

---------------------------------------------------------------
--                  Behavior Section                         --
---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);
    WBdlyd      <= WBint after 1 ps;


    PROCESS
    BEGIN
       INIT_MEM <= '1';
       WAIT;
    END PROCESS;

    VITALBehavior : process (INIT_MEM, 
                          RADDR0_ipd, RADDR1_ipd, RADDR2_ipd, RADDR3_ipd, RADDR4_ipd, RADDR5_ipd, RADDR6_ipd, RADDR7_ipd, 
                          WADDR0_ipd, WADDR1_ipd, WADDR2_ipd, WADDR3_ipd, WADDR4_ipd, WADDR5_ipd, WADDR6_ipd, WADDR7_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd 
                          )

    -- some internal veriable declaration
     variable RAM_di_int         : std_logic_vector(8 downto 0);
     variable memory_array       : MEM_TYPE := (others =>(others => 'X'));
     variable do_par             : std_logic:= 'X';
     variable tmp_par            : std_logic:= 'X';
     variable tmp_par2           : std_logic:= 'X';
     variable wpe_var            : std_logic:= 'X';

     --  Read Timing Check Results
     variable PeriodData_RDB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RDB                  : X01                 := '0';
     variable PeriodData_RBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RBLKB                : X01                  := '0';
     variable PeriodData_RADDR0          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR0               : X01                 := '0';
     variable PeriodData_RADDR1          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR1               : X01                 := '0';
     variable PeriodData_RADDR2          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR2               : X01                 := '0';
     variable PeriodData_RADDR3          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR3               : X01                 := '0';
     variable PeriodData_RADDR4          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR4               : X01                 := '0';
     variable PeriodData_RADDR5          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR5               : X01                 := '0';
     variable PeriodData_RADDR6          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR6               : X01                 := '0';
     variable PeriodData_RADDR7          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR7               : X01                 := '0';
     variable Tviol_WADDR0_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR0_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR0_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR0_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR0_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR1_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR1_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR1_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR1_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR2_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR2_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR2_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR2_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR3_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR3_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR3_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR3_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR4_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR4_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR4_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR4_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR5_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR5_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR5_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR5_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR6_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR6_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR6_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR6_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR7_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR7_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR7_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR7_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WRB_posedge      : X01                 := '0';
     variable TmDt_DI0_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI0_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WRB_posedge      : X01                 := '0';
     variable TmDt_DI1_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI1_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WRB_posedge      : X01                 := '0';
     variable TmDt_DI2_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI2_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WRB_posedge      : X01                 := '0';
     variable TmDt_DI3_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI3_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WRB_posedge      : X01                 := '0';
     variable TmDt_DI4_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI4_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WRB_posedge      : X01                 := '0';
     variable TmDt_DI5_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI5_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WRB_posedge      : X01                 := '0';
     variable TmDt_DI6_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI6_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WRB_posedge      : X01                 := '0';
     variable TmDt_DI7_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI7_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WRB_posedge      : X01                 := '0';
     variable TmDt_DI8_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI8_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WRB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WRB                  : X01                 := '0';
     variable PeriodData_WBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WBLKB                : X01                 := '0';
     variable Tviol_RDB_WRB_posedge      : X01                 := '0';
     variable TmDt_RDB_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_WRB_negedge      : X01                 := '0';
     variable TmDt_RDB_WRB_negedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_WRB_posedge    : X01                 := '0';
     variable TmDt_RBLKB_WRB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_WRB_negedge    : X01                 := '0';
     variable TmDt_RBLKB_WRB_negedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR0_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR0_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR0_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR0_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR1_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR1_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR2_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR2_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR3_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR3_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR4_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR4_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR5_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR5_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR6_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR6_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR7_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR7_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_WBLKB_posedge    : X01                 := '0';
     variable TmDt_RDB_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_WBLKB_negedge    : X01                 := '0';
     variable TmDt_RDB_WBLKB_negedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_WBLKB_posedge  : X01                 := '0';
     variable TmDt_RBLKB_WBLKB_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_WBLKB_negedge  : X01                 := '0';
     variable TmDt_RBLKB_WBLKB_negedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR0_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR0_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR0_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR0_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR1_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR1_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR2_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR2_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR3_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR3_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR4_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR4_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR5_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR5_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR6_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR6_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR7_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR7_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results

     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     variable DO0_zd : std_ulogic;
     variable DO1_zd : std_ulogic;
     variable DO2_zd : std_ulogic;
     variable DO3_zd : std_ulogic;
     variable DO4_zd : std_ulogic;
     variable DO5_zd : std_ulogic;
     variable DO6_zd : std_ulogic;
     variable DO7_zd : std_ulogic;
     variable DO8_zd : std_ulogic;
     variable RPE_zd : std_ulogic;
     variable WPE_zd : std_ulogic;
     variable DOS_zd : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData  : VitalGlitchDataType;
     variable DO1_GlitchData  : VitalGlitchDataType;
     variable DO2_GlitchData  : VitalGlitchDataType;
     variable DO3_GlitchData  : VitalGlitchDataType;
     variable DO4_GlitchData  : VitalGlitchDataType;
     variable DO5_GlitchData  : VitalGlitchDataType;
     variable DO6_GlitchData  : VitalGlitchDataType;
     variable DO7_GlitchData  : VitalGlitchDataType;
     variable DO8_GlitchData  : VitalGlitchDataType;
     variable RPE_GlitchData  : VitalGlitchDataType;
     variable WPE_GlitchData  : VitalGlitchDataType;
     variable DOS_GlitchData  : VitalGlitchDataType;

     -- last value variables
     variable RBint_previous  : std_ulogic := 'X';
     variable WBint_previous  : std_ulogic := 'X';
     variable DIS_previous    : std_ulogic := 'X';
     variable RADDR0_previous : std_ulogic := 'X';
     variable RADDR1_previous : std_ulogic := 'X';
     variable RADDR2_previous : std_ulogic := 'X';
     variable RADDR3_previous : std_ulogic := 'X';
     variable RADDR4_previous : std_ulogic := 'X';
     variable RADDR5_previous : std_ulogic := 'X';
     variable RADDR6_previous : std_ulogic := 'X';
     variable RADDR7_previous : std_ulogic := 'X';
     variable WADDR0_previous : std_ulogic := 'X';
     variable WADDR1_previous : std_ulogic := 'X';
     variable WADDR2_previous : std_ulogic := 'X';
     variable WADDR3_previous : std_ulogic := 'X';
     variable WADDR4_previous : std_ulogic := 'X';
     variable WADDR5_previous : std_ulogic := 'X';
     variable WADDR6_previous : std_ulogic := 'X';
     variable WADDR7_previous : std_ulogic := 'X';

     variable PARODD_previous : std_ulogic := 'X';
     variable Write_OK        : Boolean := FALSE;

     variable inline    : LINE;
     variable indata    : std_logic_vector(8 downto 0);
     variable resdata   : std_logic_vector(8 downto 0);
     variable i         : integer:=0;
     file     memfile   : text;
     variable status         : file_open_status;

 begin -- process VITALBehavior

  -----------------------------------------------------------
  --    Initialize memory file from MEMORYFILE string      --
  -----------------------------------------------------------

  if ( INIT_MEM'EVENT and INIT_MEM = '1') then
    file_open(status, memfile, MEMORYFILE, read_mode);
    if ( status=open_ok ) then
      while((i < 256) and (not ENDFILE(memfile))) loop
        readline(memfile,inline);
        read(inline,indata);
        resdata := indata;
        memory_array(i) := resdata;
        i := i+1;
      end loop;
    else
      assert ( MEMORYFILE'length = 0 )  
        report "Failed to open RAM256x9AA memory initialization file in read mode"
        severity Note;
    end if;
    file_close(memfile);
  end if;


      WADDR := ((INT(WADDR7_ipd)*128)+(INT(WADDR6_ipd)*64)+(INT(
               WADDR5_ipd)*32) + (INT(WADDR4_ipd)*16) + 
               (INT(WADDR3_ipd)*8) + (INT(WADDR2_ipd)*4) + (INT(
               WADDR1_ipd)*2) + (INT(WADDR0_ipd)*1));
   -- Convert Read Address Signal to Integer

      RADDR := ((INT(RADDR7_ipd)*128)+(INT(RADDR6_ipd)*64)+(INT(
               RADDR5_ipd)*32) + (INT(RADDR4_ipd)*16) + 
               (INT(RADDR3_ipd)*8) + (INT(RADDR2_ipd)*4) + (INT(
               RADDR1_ipd)*2) + (INT(RADDR0_ipd)*1));

   if ( TimingCheckOn ) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

      VitalPeriodPulseCheck ( Pviol_RDB,
                              PeriodData_RDB,
                              RDB_ipd, "RDB",
                              0.0 ns,
                              tperiod_RDB,
                              tpw_RDB_posedge,
                              tpw_RDB_negedge,
                              (To_X01(RBLKB_ipd) = '0'),
                             InstancePath &"/RAM256x9AA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RBLKB,
                              PeriodData_RBLKB,
                              RBLKB_ipd, "RBLKB",
                              0.0 ns,
                              tperiod_RBLKB,
                              tpw_RBLKB_posedge,
                              tpw_RBLKB_negedge,
                              (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR0,
                              PeriodData_RADDR0,
                              RADDR0_ipd, "RADDR0",
                              0.0 ns,
                              tpw_RADDR0_posedge + tpw_RADDR0_posedge,
                              tpw_RADDR0_posedge,
                              tpw_RADDR0_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR1,
                              PeriodData_RADDR1,
                              RADDR1_ipd, "RADDR1",
                              0.0 ns,
                              tpw_RADDR1_posedge + tpw_RADDR1_posedge,
                              tpw_RADDR1_posedge,
                              tpw_RADDR1_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR2,
                              PeriodData_RADDR2,
                              RADDR2_ipd, "RADDR2",
                              0.0 ns,
                              tpw_RADDR2_posedge + tpw_RADDR2_posedge,
                              tpw_RADDR2_posedge,
                              tpw_RADDR2_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR3,
                              PeriodData_RADDR3,
                              RADDR3_ipd, "RADDR3",
                              0.0 ns,
                              tpw_RADDR3_posedge + tpw_RADDR3_posedge,
                              tpw_RADDR3_posedge,
                              tpw_RADDR3_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR4,
                              PeriodData_RADDR4,
                              RADDR4_ipd, "RADDR4",
                              0.0 ns,
                              tpw_RADDR4_posedge + tpw_RADDR4_posedge,
                              tpw_RADDR4_posedge,
                              tpw_RADDR4_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR5,
                              PeriodData_RADDR5,
                              RADDR5_ipd, "RADDR5",
                              0.0 ns,
                              tpw_RADDR5_posedge + tpw_RADDR5_posedge,
                              tpw_RADDR5_posedge,
                              tpw_RADDR5_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR6,
                              PeriodData_RADDR6,
                              RADDR6_ipd, "RADDR6",
                              0.0 ns,
                              tpw_RADDR6_posedge + tpw_RADDR6_posedge,
                              tpw_RADDR6_posedge,
                              tpw_RADDR6_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR7,
                              PeriodData_RADDR7,
                              RADDR7_ipd, "RADDR7",
                              0.0 ns,
                              tpw_RADDR7_posedge + tpw_RADDR7_posedge,
                              tpw_RADDR7_posedge,
                              tpw_RADDR7_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AA",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_negedge,
                             TmDt_WADDR0_WRB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR0_WRB_posedge_negedge,
                             tsetup_WADDR0_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_negedge,
                             TmDt_WADDR0_WRB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR0_WRB_negedge_negedge,
                             tsetup_WADDR0_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_negedge,
                             TmDt_WADDR1_WRB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR1_WRB_posedge_negedge,
                             tsetup_WADDR1_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_negedge,
                             TmDt_WADDR1_WRB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR1_WRB_negedge_negedge,
                             tsetup_WADDR1_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_negedge,
                             TmDt_WADDR2_WRB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR2_WRB_posedge_negedge,
                             tsetup_WADDR2_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_negedge,
                             TmDt_WADDR2_WRB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR2_WRB_negedge_negedge,
                             tsetup_WADDR2_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_negedge,
                             TmDt_WADDR3_WRB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR3_WRB_posedge_negedge,
                             tsetup_WADDR3_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_negedge,
                             TmDt_WADDR3_WRB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR3_WRB_negedge_negedge,
                             tsetup_WADDR3_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_negedge,
                             TmDt_WADDR4_WRB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR4_WRB_posedge_negedge,
                             tsetup_WADDR4_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_negedge,
                             TmDt_WADDR4_WRB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR4_WRB_negedge_negedge,
                             tsetup_WADDR4_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_negedge,
                             TmDt_WADDR5_WRB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR5_WRB_posedge_negedge,
                             tsetup_WADDR5_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_negedge,
                             TmDt_WADDR5_WRB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR5_WRB_negedge_negedge,
                             tsetup_WADDR5_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_negedge,
                             TmDt_WADDR6_WRB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR6_WRB_posedge_negedge,
                             tsetup_WADDR6_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_negedge,
                             TmDt_WADDR6_WRB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR6_WRB_negedge_negedge,
                             tsetup_WADDR6_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_negedge,
                             TmDt_WADDR7_WRB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR7_WRB_posedge_negedge,
                             tsetup_WADDR7_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_negedge,
                             TmDt_WADDR7_WRB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR7_WRB_negedge_negedge,
                             tsetup_WADDR7_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_negedge,
                             TmDt_WADDR0_WBLKB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR0_WBLKB_posedge_negedge,
                             tsetup_WADDR0_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_negedge,
                             TmDt_WADDR0_WBLKB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR0_WBLKB_negedge_negedge,
                             tsetup_WADDR0_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_negedge,
                             TmDt_WADDR1_WBLKB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR1_WBLKB_posedge_negedge,
                             tsetup_WADDR1_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_negedge,
                             TmDt_WADDR1_WBLKB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR1_WBLKB_negedge_negedge,
                             tsetup_WADDR1_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_negedge,
                             TmDt_WADDR2_WBLKB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR2_WBLKB_posedge_negedge,
                             tsetup_WADDR2_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_negedge,
                             TmDt_WADDR2_WBLKB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR2_WBLKB_negedge_negedge,
                             tsetup_WADDR2_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_negedge,
                             TmDt_WADDR3_WBLKB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR3_WBLKB_posedge_negedge,
                             tsetup_WADDR3_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_negedge,
                             TmDt_WADDR3_WBLKB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR3_WBLKB_negedge_negedge,
                             tsetup_WADDR3_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_negedge,
                             TmDt_WADDR4_WBLKB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR4_WBLKB_posedge_negedge,
                             tsetup_WADDR4_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_negedge,
                             TmDt_WADDR4_WBLKB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR4_WBLKB_negedge_negedge,
                             tsetup_WADDR4_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_negedge,
                             TmDt_WADDR5_WBLKB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR5_WBLKB_posedge_negedge,
                             tsetup_WADDR5_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_negedge,
                             TmDt_WADDR5_WBLKB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR5_WBLKB_negedge_negedge,
                             tsetup_WADDR5_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_negedge,
                             TmDt_WADDR6_WBLKB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR6_WBLKB_posedge_negedge,
                             tsetup_WADDR6_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_negedge,
                             TmDt_WADDR6_WBLKB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR6_WBLKB_negedge_negedge,
                             tsetup_WADDR6_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_negedge,
                             TmDt_WADDR7_WBLKB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR7_WBLKB_posedge_negedge,
                             tsetup_WADDR7_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_negedge,
                             TmDt_WADDR7_WBLKB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR7_WBLKB_negedge_negedge,
                             tsetup_WADDR7_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_posedge,
                             TmDt_WADDR0_WRB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WRB_posedge_posedge,
                             thold_WADDR0_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_posedge,
                             TmDt_WADDR0_WRB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WRB_negedge_posedge,
                             thold_WADDR0_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_posedge,
                             TmDt_WADDR1_WRB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WRB_posedge_posedge,
                             thold_WADDR1_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_posedge,
                             TmDt_WADDR1_WRB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WRB_negedge_posedge,
                             thold_WADDR1_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_posedge,
                             TmDt_WADDR2_WRB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WRB_posedge_posedge,
                             thold_WADDR2_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_posedge,
                             TmDt_WADDR2_WRB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WRB_negedge_posedge,
                             thold_WADDR2_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_posedge,
                             TmDt_WADDR3_WRB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WRB_posedge_posedge,
                             thold_WADDR3_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_posedge,
                             TmDt_WADDR3_WRB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WRB_negedge_posedge,
                             thold_WADDR3_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_posedge,
                             TmDt_WADDR4_WRB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WRB_posedge_posedge,
                             thold_WADDR4_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_posedge,
                             TmDt_WADDR4_WRB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WRB_negedge_posedge,
                             thold_WADDR4_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_posedge,
                             TmDt_WADDR5_WRB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WRB_posedge_posedge,
                             thold_WADDR5_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_posedge,
                             TmDt_WADDR5_WRB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WRB_negedge_posedge,
                             thold_WADDR5_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_posedge,
                             TmDt_WADDR6_WRB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WRB_posedge_posedge,
                             thold_WADDR6_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_posedge,
                             TmDt_WADDR6_WRB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WRB_negedge_posedge,
                             thold_WADDR6_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_posedge,
                             TmDt_WADDR7_WRB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WRB_posedge_posedge,
                             thold_WADDR7_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_posedge,
                             TmDt_WADDR7_WRB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WRB_negedge_posedge,
                             thold_WADDR7_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_posedge,
                             TmDt_WADDR0_WBLKB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WBLKB_posedge_posedge,
                             thold_WADDR0_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_posedge,
                             TmDt_WADDR0_WBLKB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WBLKB_negedge_posedge,
                             thold_WADDR0_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_posedge,
                             TmDt_WADDR1_WBLKB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WBLKB_posedge_posedge,
                             thold_WADDR1_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_posedge,
                             TmDt_WADDR1_WBLKB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WBLKB_negedge_posedge,
                             thold_WADDR1_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_posedge,
                             TmDt_WADDR2_WBLKB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WBLKB_posedge_posedge,
                             thold_WADDR2_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_posedge,
                             TmDt_WADDR2_WBLKB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WBLKB_negedge_posedge,
                             thold_WADDR2_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_posedge,
                             TmDt_WADDR3_WBLKB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WBLKB_posedge_posedge,
                             thold_WADDR3_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_posedge,
                             TmDt_WADDR3_WBLKB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WBLKB_negedge_posedge,
                             thold_WADDR3_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_posedge,
                             TmDt_WADDR4_WBLKB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WBLKB_posedge_posedge,
                             thold_WADDR4_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_posedge,
                             TmDt_WADDR4_WBLKB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WBLKB_negedge_posedge,
                             thold_WADDR4_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_posedge,
                             TmDt_WADDR5_WBLKB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WBLKB_posedge_posedge,
                             thold_WADDR5_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_posedge,
                             TmDt_WADDR5_WBLKB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WBLKB_negedge_posedge,
                             thold_WADDR5_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_posedge,
                             TmDt_WADDR6_WBLKB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WBLKB_posedge_posedge,
                             thold_WADDR6_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_posedge,
                             TmDt_WADDR6_WBLKB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WBLKB_negedge_posedge,
                             thold_WADDR6_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_posedge,
                             TmDt_WADDR7_WBLKB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WBLKB_posedge_posedge,
                             thold_WADDR7_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_posedge,
                             TmDt_WADDR7_WBLKB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WBLKB_negedge_posedge,
                             thold_WADDR7_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_posedge_posedge,
                             tsetup_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_negedge_posedge,
                             tsetup_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_posedge_posedge,
                             tsetup_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_negedge_posedge,
                             tsetup_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_posedge_posedge,
                             tsetup_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_negedge_posedge,
                             tsetup_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_posedge_posedge,
                             tsetup_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_negedge_posedge,
                             tsetup_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_posedge_posedge,
                             tsetup_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_negedge_posedge,
                             tsetup_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_posedge_posedge,
                             tsetup_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_negedge_posedge,
                             tsetup_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_posedge_posedge,
                             tsetup_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_negedge_posedge,
                             tsetup_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_posedge_posedge,
                             tsetup_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_negedge_posedge,
                             tsetup_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_posedge_posedge,
                             tsetup_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_negedge_posedge,
                             tsetup_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_posedge_posedge,
                             tsetup_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_negedge_posedge,
                             tsetup_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_posedge_posedge,
                             tsetup_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_negedge_posedge,
                             tsetup_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_posedge_posedge,
                             tsetup_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_negedge_posedge,
                             tsetup_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_posedge_posedge,
                             tsetup_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_negedge_posedge,
                             tsetup_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_posedge_posedge,
                             tsetup_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_negedge_posedge,
                             tsetup_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_posedge_posedge,
                             tsetup_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_negedge_posedge,
                             tsetup_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_posedge_posedge,
                             tsetup_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_negedge_posedge,
                             tsetup_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_posedge_posedge,
                             tsetup_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_negedge_posedge,
                             tsetup_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_posedge_posedge,
                             tsetup_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_negedge_posedge,
                             tsetup_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AA",
                             True,
                             True,
                             WARNING
                             );
      VitalPeriodPulseCheck ( Pviol_WBLKB,
                              PeriodData_WBLKB,
                              WBLKB_ipd, "WBLKB",
                              0.0 ns,
                              tperiod_WBLKB,
                              tpw_WBLKB_posedge,
                              tpw_WBLKB_negedge,
                              (To_X01(WRB_ipd) = '0'),
                              InstancePath & "/RAM256x9AA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_WRB,
                              PeriodData_WRB,
                              WRB_ipd, "WRB",
                              0.0 ns,
                              tperiod_WRB,
                              tpw_WRB_posedge,
                              tpw_WRB_negedge,
                              (To_X01(WBLKB_ipd) = '0'),
                              InstancePath & "/RAM256x9AA",
                              True,
                              True,
                              WARNING
                              );
   ------------------------------------------------------------
   --        Timing Checking for Read and write conflict     --
   ------------------------------------------------------------
       VitalSetupHoldCheck ( Tviol_RDB_WRB_negedge,
                             TmDt_RDB_WRB_negedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_RDB_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_WBLKB_negedge,
                             TmDt_RDB_WBLKB_negedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_RDB_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB) = '0') AND (To_X01(RBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_WRB_posedge,
                             TmDt_RDB_WRB_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RDB_WRB_posedge_posedge,
                             0.0 ns,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_WBLKB_posedge,
                             TmDt_RDB_WBLKB_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RDB_WBLKB_posedge_posedge,
                             0.0 ns,
                             (To_X01(WRB) = '0') AND (To_X01(RBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_WRB_negedge,
                             TmDt_RBLKB_WRB_negedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_RBLKB_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB) = '0') AND (To_X01(RDB_ipd) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_WBLKB_negedge,
                             TmDt_RBLKB_WBLKB_negedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_RBLKB_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB) = '0') AND (To_X01(RDB_ipd) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_WRB_posedge,
                             TmDt_RBLKB_WRB_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RBLKB_WRB_posedge_posedge,
                             0.0 ns,
                             (To_X01(WBLKB) = '0') AND (To_X01(RDB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_WBLKB_posedge,
                             TmDt_RBLKB_WBLKB_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RBLKB_WBLKB_posedge_posedge,
                             0.0 ns,
                             (To_X01(WRB) = '0') AND (To_X01(RDB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WRB_posedge,
                             TmDt_RADDR0_WRB_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR0_WRB_negedge_posedge,
                             thold_RADDR0_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WRB_posedge,
                             TmDt_RADDR0_WRB_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR0_WRB_posedge_posedge,
                             thold_RADDR0_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WRB_negedge,
                             TmDt_RADDR0_WRB_negedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR0_WRB_posedge_negedge,
                             tsetup_RADDR0_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WRB_negedge,
                             TmDt_RADDR0_WRB_negedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR0_WRB_negedge_negedge,
                             tsetup_RADDR0_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WBLKB_posedge,
                             TmDt_RADDR0_WBLKB_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR0_WRB_negedge_posedge,
                             thold_RADDR0_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WBLKB_posedge,
                             TmDt_RADDR0_WBLKB_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR0_WRB_posedge_posedge,
                             thold_RADDR0_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WBLKB_negedge,
                             TmDt_RADDR0_WBLKB_negedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR0_WBLKB_posedge_negedge,
                             tsetup_RADDR0_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WBLKB_negedge,
                             TmDt_RADDR0_WBLKB_negedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR0_WBLKB_negedge_negedge,
                             tsetup_RADDR0_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WRB_posedge,
                             TmDt_RADDR1_WRB_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR1_WRB_negedge_posedge,
                             thold_RADDR1_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WRB_posedge,
                             TmDt_RADDR1_WRB_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR1_WRB_posedge_posedge,
                             thold_RADDR1_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WRB_negedge,
                             TmDt_RADDR1_WRB_negedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR1_WRB_posedge_negedge,
                             tsetup_RADDR1_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WRB_negedge,
                             TmDt_RADDR1_WRB_negedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR1_WRB_negedge_negedge,
                             tsetup_RADDR1_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WBLKB_posedge,
                             TmDt_RADDR1_WBLKB_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR1_WRB_negedge_posedge,
                             thold_RADDR1_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WBLKB_posedge,
                             TmDt_RADDR1_WBLKB_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR1_WRB_posedge_posedge,
                             thold_RADDR1_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WBLKB_negedge,
                             TmDt_RADDR1_WBLKB_negedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR1_WBLKB_posedge_negedge,
                             tsetup_RADDR1_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WBLKB_negedge,
                             TmDt_RADDR1_WBLKB_negedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR1_WBLKB_negedge_negedge,
                             tsetup_RADDR1_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WRB_posedge,
                             TmDt_RADDR2_WRB_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR2_WRB_negedge_posedge,
                             thold_RADDR2_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WRB_posedge,
                             TmDt_RADDR2_WRB_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR2_WRB_posedge_posedge,
                             thold_RADDR2_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WRB_negedge,
                             TmDt_RADDR2_WRB_negedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR2_WRB_posedge_negedge,
                             tsetup_RADDR2_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WRB_negedge,
                             TmDt_RADDR2_WRB_negedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR2_WRB_negedge_negedge,
                             tsetup_RADDR2_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WBLKB_posedge,
                             TmDt_RADDR2_WBLKB_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR2_WRB_negedge_posedge,
                             thold_RADDR2_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WBLKB_posedge,
                             TmDt_RADDR2_WBLKB_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR2_WRB_posedge_posedge,
                             thold_RADDR2_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WBLKB_negedge,
                             TmDt_RADDR2_WBLKB_negedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR2_WBLKB_posedge_negedge,
                             tsetup_RADDR2_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WBLKB_negedge,
                             TmDt_RADDR2_WBLKB_negedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR2_WBLKB_negedge_negedge,
                             tsetup_RADDR2_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WRB_posedge,
                             TmDt_RADDR3_WRB_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR3_WRB_negedge_posedge,
                             thold_RADDR3_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WRB_posedge,
                             TmDt_RADDR3_WRB_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR3_WRB_posedge_posedge,
                             thold_RADDR3_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WRB_negedge,
                             TmDt_RADDR3_WRB_negedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR3_WRB_posedge_negedge,
                             tsetup_RADDR3_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WRB_negedge,
                             TmDt_RADDR3_WRB_negedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR3_WRB_negedge_negedge,
                             tsetup_RADDR3_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WBLKB_posedge,
                             TmDt_RADDR3_WBLKB_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR3_WRB_negedge_posedge,
                             thold_RADDR3_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WBLKB_posedge,
                             TmDt_RADDR3_WBLKB_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR3_WRB_posedge_posedge,
                             thold_RADDR3_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WBLKB_negedge,
                             TmDt_RADDR3_WBLKB_negedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR3_WBLKB_posedge_negedge,
                             tsetup_RADDR3_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WBLKB_negedge,
                             TmDt_RADDR3_WBLKB_negedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR3_WBLKB_negedge_negedge,
                             tsetup_RADDR3_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WRB_posedge,
                             TmDt_RADDR4_WRB_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR4_WRB_negedge_posedge,
                             thold_RADDR4_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WRB_posedge,
                             TmDt_RADDR4_WRB_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR4_WRB_posedge_posedge,
                             thold_RADDR4_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WRB_negedge,
                             TmDt_RADDR4_WRB_negedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR4_WRB_posedge_negedge,
                             tsetup_RADDR4_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WRB_negedge,
                             TmDt_RADDR4_WRB_negedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR4_WRB_negedge_negedge,
                             tsetup_RADDR4_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WBLKB_posedge,
                             TmDt_RADDR4_WBLKB_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR4_WRB_negedge_posedge,
                             thold_RADDR4_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WBLKB_posedge,
                             TmDt_RADDR4_WBLKB_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR4_WRB_posedge_posedge,
                             thold_RADDR4_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WBLKB_negedge,
                             TmDt_RADDR4_WBLKB_negedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR4_WBLKB_posedge_negedge,
                             tsetup_RADDR4_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WBLKB_negedge,
                             TmDt_RADDR4_WBLKB_negedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR4_WBLKB_negedge_negedge,
                             tsetup_RADDR4_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WRB_posedge,
                             TmDt_RADDR5_WRB_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR5_WRB_negedge_posedge,
                             thold_RADDR5_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WRB_posedge,
                             TmDt_RADDR5_WRB_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR5_WRB_posedge_posedge,
                             thold_RADDR5_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WRB_negedge,
                             TmDt_RADDR5_WRB_negedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR5_WRB_posedge_negedge,
                             tsetup_RADDR5_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WRB_negedge,
                             TmDt_RADDR5_WRB_negedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR5_WRB_negedge_negedge,
                             tsetup_RADDR5_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WBLKB_posedge,
                             TmDt_RADDR5_WBLKB_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR5_WRB_negedge_posedge,
                             thold_RADDR5_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WBLKB_posedge,
                             TmDt_RADDR5_WBLKB_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR5_WRB_posedge_posedge,
                             thold_RADDR5_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WBLKB_negedge,
                             TmDt_RADDR5_WBLKB_negedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR5_WBLKB_posedge_negedge,
                             tsetup_RADDR5_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WBLKB_negedge,
                             TmDt_RADDR5_WBLKB_negedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR5_WBLKB_negedge_negedge,
                             tsetup_RADDR5_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WRB_posedge,
                             TmDt_RADDR6_WRB_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR6_WRB_negedge_posedge,
                             thold_RADDR6_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WRB_posedge,
                             TmDt_RADDR6_WRB_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR6_WRB_posedge_posedge,
                             thold_RADDR6_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WRB_negedge,
                             TmDt_RADDR6_WRB_negedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR6_WRB_posedge_negedge,
                             tsetup_RADDR6_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WRB_negedge,
                             TmDt_RADDR6_WRB_negedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR6_WRB_negedge_negedge,
                             tsetup_RADDR6_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WBLKB_posedge,
                             TmDt_RADDR6_WBLKB_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR6_WRB_negedge_posedge,
                             thold_RADDR6_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WBLKB_posedge,
                             TmDt_RADDR6_WBLKB_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR6_WRB_posedge_posedge,
                             thold_RADDR6_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WBLKB_negedge,
                             TmDt_RADDR6_WBLKB_negedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR6_WBLKB_posedge_negedge,
                             tsetup_RADDR6_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WBLKB_negedge,
                             TmDt_RADDR6_WBLKB_negedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR6_WBLKB_negedge_negedge,
                             tsetup_RADDR6_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WRB_posedge,
                             TmDt_RADDR7_WRB_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR7_WRB_negedge_posedge,
                             thold_RADDR7_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WRB_posedge,
                             TmDt_RADDR7_WRB_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR7_WRB_posedge_posedge,
                             thold_RADDR7_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WRB_negedge,
                             TmDt_RADDR7_WRB_negedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR7_WRB_posedge_negedge,
                             tsetup_RADDR7_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WRB_negedge,
                             TmDt_RADDR7_WRB_negedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR7_WRB_negedge_negedge,
                             tsetup_RADDR7_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WBLKB_posedge,
                             TmDt_RADDR7_WBLKB_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR7_WRB_negedge_posedge,
                             thold_RADDR7_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WBLKB_posedge,
                             TmDt_RADDR7_WBLKB_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR7_WRB_posedge_posedge,
                             thold_RADDR7_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WBLKB_negedge,
                             TmDt_RADDR7_WBLKB_negedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR7_WBLKB_posedge_negedge,
                             tsetup_RADDR7_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WBLKB_negedge,
                             TmDt_RADDR7_WBLKB_negedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR7_WBLKB_negedge_negedge,
                             tsetup_RADDR7_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

   end if;

   ------------------------------------------------------------
   --    wpe output                                           -
   ------------------------------------------------------------

   if ( PARODD_ipd'EVENT ) then
     RPE_zd := not RPE_zd;
     WPE_zd := not WPE_zd;
   end if;

   ------------------------------------------------------------
   --         WPE checking  block                            -
   ------------------------------------------------------------

      tmp_par  := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;
      tmp_par2 := (tmp_par xor DI8_ipd);

      if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
          ( TO_X01 ( DI8_ipd )    = 'X' ) or
          ( TO_X01 ( DI7_ipd )    = 'X' ) or
          ( TO_X01 ( DI6_ipd )    = 'X' ) or
          ( TO_X01 ( DI5_ipd )    = 'X' ) or
          ( TO_X01 ( DI4_ipd )    = 'X' ) or
          ( TO_X01 ( DI3_ipd )    = 'X' ) or
          ( TO_X01 ( DI2_ipd )    = 'X' ) or
          ( TO_X01 ( DI1_ipd )    = 'X' ) or
          ( TO_X01 ( DI0_ipd )    = 'X' )
         ) then
        wpe_var  :=  'X';
      else
        if ( tmp_par2 /= PARODD_ipd ) then
          wpe_var  :=  '1';
        else
          wpe_var  :=  '0';
        end if;
      end if;
      RAM_di_int(8) := DI8_ipd;
      WPE_zd := wpe_var;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

    if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
    end if; 

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------
   
   if (( TO_X01 ( WBint ) = '0' ) and ( TO_X01 ( WBint_previous ) = '1' )) then
     Write_OK := True;
   end if;

 -- async memory writing 
   if ( WBint'event or WADDR0_ipd'event or WADDR1_ipd'event or 
        WADDR2_ipd'event or WADDR3_ipd'event or WADDR4_ipd'event or 
        WADDR5_ipd'event or WADDR6_ipd'event or WADDR7_ipd'event or 
        DI7_ipd'event or DI6_ipd'event or DI5_ipd'event or 
        DI4_ipd'event or DI3_ipd'event or DI2_ipd'event or 
        DI1_ipd'event or DI0_ipd'event or DI8_ipd'event ) then
     if (TO_X01(WBint)='X') then
       if (TO_X01(WBint_previous) /= 'X') then
         assert false
           report ": WRB or WBLKB unknown"
           severity Warning;
       end if;
     elsif ( TO_X01(WBint) = '0' and Write_OK ) then
       if(WADDR < 0) then
           if((TO_X01(WADDR0_ipd) = 'X') and (TO_X01(WADDR0_previous) /= 'X')) then
             assert false
             report ": WADDR0 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR1_ipd) = 'X') and (TO_X01(WADDR1_previous) /= 'X')) then
             assert false
             report ": WADDR1 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR2_ipd) = 'X') and (TO_X01(WADDR2_previous) /= 'X')) then
             assert false
             report ": WADDR2 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR3_ipd) = 'X') and (TO_X01(WADDR3_previous) /= 'X')) then
             assert false
             report ": WADDR3 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR4_ipd) = 'X') and (TO_X01(WADDR4_previous) /= 'X')) then
             assert false
             report ": WADDR4 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR5_ipd) = 'X') and (TO_X01(WADDR5_previous) /= 'X')) then
             assert false
             report ": WADDR5 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR6_ipd) = 'X') and (TO_X01(WADDR6_previous) /= 'X')) then
             assert false
             report ": WADDR6 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR7_ipd) = 'X') and (TO_X01(WADDR7_previous) /= 'X')) then
             assert false
             report ": WADDR7 unknown, no data written ......"
             severity Warning;
           end if;
       else
         RAM_di_int ( 7 downto 0 ) := DI7_ipd & DI6_ipd & DI5_ipd & DI4_ipd & 
                                      DI3_ipd & DI2_ipd & DI1_ipd & DI0_ipd;
         memory_array ( WADDR ) := RAM_di_int;
       end if;
     end if;
   end if;


 -----------------------------------------------------------
 --  Read Functional Section                              --
 -----------------------------------------------------------



-- Asynchronous RAM Read, Enable signal controlled;

   if ( RBint'event or RADDR0_ipd'event or RADDR1_ipd'event or 
        RADDR2_ipd'event or RADDR3_ipd'event or RADDR4_ipd'event or 
        RADDR5_ipd'event or RADDR6_ipd'event or RADDR7_ipd'event or
        WBint'event or WADDR0_ipd'event or WADDR1_ipd'event or 
        WADDR2_ipd'event or WADDR3_ipd'event or WADDR4_ipd'event or 
        WADDR5_ipd'event or WADDR6_ipd'event or WADDR7_ipd'event
      ) then
     if ( TO_X01 ( RBint ) = 'X' ) then
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          RPE_zd :='X';
          if ( TO_X01 ( RBint_previous ) /= 'X' ) then
             assert false
               report ": RDB or RBLKB unknown"
               severity Warning;
          end if;
     elsif ( RADDR < 0 ) then
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          RPE_zd :='X';
          if(TO_X01(RADDR0_ipd) = 'X') and (TO_X01(RADDR0_previous) /= 'X') then
             assert false
             report ": RADDR0 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR1_ipd) = 'X') and (TO_X01(RADDR1_previous) /= 'X') then
             assert false
             report ": RADDR1 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR2_ipd) = 'X') and (TO_X01(RADDR2_previous) /= 'X') then
             assert false
             report ": RADDR2 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR3_ipd) = 'X') and (TO_X01(RADDR3_previous) /= 'X') then
             assert false
             report ": RADDR3 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR4_ipd) = 'X') and (TO_X01(RADDR4_previous) /= 'X') then
             assert false
             report ": RADDR4 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR5_ipd) = 'X') and (TO_X01(RADDR5_previous) /= 'X') then
             assert false
             report ": RADDR5 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR6_ipd) = 'X') and (TO_X01(RADDR6_previous) /= 'X') then
             assert false
             report ": RADDR6 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR7_ipd) = 'X') and (TO_X01(RADDR7_previous) /= 'X') then
             assert false
             report ": RADDR7 unknown"
             severity Warning;
          end if;
     elsif ( WADDR = RADDR ) then
       if (( RBint'event AND ( TO_X01 ( RBint ) = '0' ) AND ( TO_X01 ( WBint ) = '1' )) OR
           ( WBint'event AND ( TO_X01 ( WBint ) = '1' ) AND ( TO_X01 ( RBint ) = '0' )) OR
           --( RBint'event AND ( TO_X01 ( RBint ) = '1' ) AND ( TO_X01 ( WBint ) = '0' )) OR
           ( RBint'event AND ( TO_X01 ( RBint ) = '1' ) AND ( TO_X01 ( WBdlyd ) = '0' )) OR
           (( TO_X01 ( WBint ) = '1' ) AND ( TO_X01 ( RBint ) = '0' ) AND 
            ( RADDR0_ipd'event or RADDR1_ipd'event or 
              RADDR2_ipd'event or RADDR3_ipd'event or RADDR4_ipd'event or 
              RADDR5_ipd'event or RADDR6_ipd'event or RADDR7_ipd'event ))
          ) then
             DO0_zd := memory_array(RADDR)(0);
             DO1_zd := memory_array(RADDR)(1);
             DO2_zd := memory_array(RADDR)(2);
             DO3_zd := memory_array(RADDR)(3);
             DO4_zd := memory_array(RADDR)(4);
             DO5_zd := memory_array(RADDR)(5);
             DO6_zd := memory_array(RADDR)(6);
             DO7_zd := memory_array(RADDR)(7);
             DO8_zd := memory_array(RADDR)(8);
             do_par := DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR 
                       DO3_zd XOR DO2_zd XOR DO1_zd XOR DO0_zd;
             if (do_par = 'X') then
               RPE_zd := 'X';
             elsif (do_par /= PARODD_ipd) then
               RPE_zd := '1';
             else
               RPE_zd :=  '0';
             end if;
       end if;
     else -- WADDR /= RADDR
       if ((( TO_X01 ( WBint ) = '0' ) AND ( TO_X01 ( RBint ) = '0' ) AND
            ( RADDR0_ipd'event or RADDR1_ipd'event or RADDR2_ipd'event or 
              RADDR3_ipd'event or RADDR4_ipd'event or RADDR5_ipd'event or 
              RADDR6_ipd'event or RADDR7_ipd'event or WADDR0_ipd'event or 
              WADDR1_ipd'event or WADDR2_ipd'event or WADDR3_ipd'event or 
              WADDR4_ipd'event or WADDR5_ipd'event or WADDR6_ipd'event or 
              WADDR7_ipd'event)) OR
           ( RBint'event AND ( TO_X01 ( RBint ) = '0' )) OR
           (( TO_X01 ( RBint ) = '0' ) AND
            ( RADDR0_ipd'event or RADDR1_ipd'event or RADDR2_ipd'event or 
              RADDR3_ipd'event or RADDR4_ipd'event or RADDR5_ipd'event or 
              RADDR6_ipd'event or RADDR7_ipd'event or WADDR0_ipd'event or 
              WADDR1_ipd'event or WADDR2_ipd'event or WADDR3_ipd'event or 
              WADDR4_ipd'event or WADDR5_ipd'event or WADDR6_ipd'event or 
              WADDR7_ipd'event))
          ) then
             DO0_zd := memory_array(RADDR)(0);
             DO1_zd := memory_array(RADDR)(1);
             DO2_zd := memory_array(RADDR)(2);
             DO3_zd := memory_array(RADDR)(3);
             DO4_zd := memory_array(RADDR)(4);
             DO5_zd := memory_array(RADDR)(5);
             DO6_zd := memory_array(RADDR)(6);
             DO7_zd := memory_array(RADDR)(7);
             DO8_zd := memory_array(RADDR)(8);
             do_par := DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR 
                       DO3_zd XOR DO2_zd XOR DO1_zd XOR DO0_zd;
             if (do_par = 'X') then
               RPE_zd := 'X';
             elsif (do_par /= PARODD_ipd) then
               RPE_zd := '1';
             else
               RPE_zd :=  '0';
             end if;
       end if;
     end if;
   end if;


  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       RBint_previous  := RBint;
       WBint_previous  := WBint;
       RADDR0_previous := RADDR0_ipd;
       RADDR1_previous := RADDR1_ipd;
       RADDR2_previous := RADDR2_ipd;
       RADDR3_previous := RADDR3_ipd;
       RADDR4_previous := RADDR4_ipd;
       RADDR5_previous := RADDR5_ipd;
       RADDR6_previous := RADDR6_ipd;
       RADDR7_previous := RADDR7_ipd;
       WADDR0_previous := WADDR0_ipd;
       WADDR1_previous := WADDR1_ipd;
       WADDR2_previous := WADDR2_ipd;
       WADDR3_previous := WADDR3_ipd;
       WADDR4_previous := WADDR4_ipd;
       WADDR5_previous := WADDR5_ipd;
       WADDR6_previous := WADDR6_ipd;
       WADDR7_previous := WADDR7_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
           OutSignal     => DOS,
           GlitchData    => DOS_GlitchData,
           OutSignalName => "DOS",
           OutTemp       => DOS_zd,
           Paths  =>  (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),
           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => WPE,
           GlitchData    => WPE_GlitchData,
           OutSignalName => "WPE",
           OutTemp       => WPE_zd,

           Paths  =>   (0 => (DI0_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI0_WPE),true),
                        1 => (DI1_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI1_WPE), true),
                        2 => (DI2_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI2_WPE), true),
                        3 => (DI3_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI3_WPE), true),
                        4 => (DI4_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI4_WPE), true),
                        5 => (DI5_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI5_WPE), true),
                        6 => (DI6_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI6_WPE), true),
                        7 => (DI7_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI7_WPE), true),
                        8 => (DI8_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI8_WPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO0), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO0), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO0), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO0), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO0), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO0), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO0), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO0), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO0), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO1), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO1), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO1), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO1), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO1), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO1), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO1), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO1), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO1), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO2), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO2), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO2), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO2), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO2), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO2), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO2), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO2), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO2), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO3), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO3), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO3), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO3), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO3), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO3), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO3), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO3), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO3), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO4), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO4), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO4), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO4), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO4), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO4), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO4), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO4), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO4), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO5), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO5), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO5), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO5), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO5), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO5), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO5), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO5), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO5), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO6), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO6), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO6), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO6), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO6), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO6), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO6), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO6), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO6), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO7), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO7), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO7), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO7), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO7), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO7), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO7), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO7), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO7), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO8), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO8), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO8), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO8), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO8), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO8), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO8), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO8), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO8), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => RPE,
           GlitchData    => RPE_GlitchData,
           OutSignalName => "RPE",
           OutTemp       => RPE_zd,

           Paths  =>   (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_RPE), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_RPE), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_RPE), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_RPE), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_RPE), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_RPE), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_RPE), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_RPE), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_RPE), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_RPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

   end process VITALBehavior;

 end VITAL_ACT;
 
 configuration CFG_RAM256x9AA_VITAL of RAM256x9AA is
    for VITAL_ACT
    end for;
 end CFG_RAM256x9AA_VITAL;


---- CELL RAM256x9AAP ----

LIBRARY ieee;
LIBRARY STD;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

USE std.textio.all;
USE ieee.std_logic_textio.all;
LIBRARY a500k;
USE a500k.all;

entity RAM256x9AAP is 

   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpw_RDB_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_RDB_negedge	        : VitalDelayType := 0.000 ns;
 	tperiod_RDB	        : VitalDelayType := 0.000 ns;
 	tpw_RBLKB_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RBLKB_negedge	: VitalDelayType := 0.000 ns;
 	tperiod_RBLKB	        : VitalDelayType := 0.000 ns;
 	tpw_RADDR0_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR0_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                           : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                         : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                         : VitalDelayType := 0.000 ns;
 	tperiod_WRB                             : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_RDB_WRB_negedge_negedge          : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_WRB_posedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RBLKB_WRB_posedge_posedge         : VitalDelayType := 0.000 ns;
 	thold_RDB_WBLKB_posedge_posedge         : VitalDelayType := 0.000 ns;
 	thold_RBLKB_WBLKB_posedge_posedge       : VitalDelayType := 0.000 ns;
 	thold_RADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
        thold_RADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');

ATTRIBUTE VITAL_LEVEL0 OF RAM256x9AAP : entity IS True ;
END RAM256x9AAP;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of RAM256x9AAP is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal WADDR0_ipd : std_ulogic := 'X';
   signal WADDR1_ipd : std_ulogic := 'X';
   signal WADDR2_ipd : std_ulogic := 'X';
   signal WADDR3_ipd : std_ulogic := 'X';
   signal WADDR4_ipd : std_ulogic := 'X';
   signal WADDR5_ipd : std_ulogic := 'X';
   signal WADDR6_ipd : std_ulogic := 'X';
   signal WADDR7_ipd : std_ulogic := 'X';
   signal RADDR0_ipd : std_ulogic := 'X';
   signal RADDR1_ipd : std_ulogic := 'X';
   signal RADDR2_ipd : std_ulogic := 'X';
   signal RADDR3_ipd : std_ulogic := 'X';
   signal RADDR4_ipd : std_ulogic := 'X';
   signal RADDR5_ipd : std_ulogic := 'X';
   signal RADDR6_ipd : std_ulogic := 'X';
   signal RADDR7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

	-- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';
   signal INIT_MEM   : std_logic:= '0';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic:= 'X';
   signal par_f2     : std_logic:= 'X';
   signal WBdlyd     : std_ulogic := 'X';

 begin  --  VITAL_ACT
   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (WADDR0_ipd, WADDR0, VitalExtendToFillDelay(tipd_WADDR0));
   VitalWireDelay (WADDR1_ipd, WADDR1, VitalExtendToFillDelay(tipd_WADDR1));
   VitalWireDelay (WADDR2_ipd, WADDR2, VitalExtendToFillDelay(tipd_WADDR2));
   VitalWireDelay (WADDR3_ipd, WADDR3, VitalExtendToFillDelay(tipd_WADDR3));
   VitalWireDelay (WADDR4_ipd, WADDR4, VitalExtendToFillDelay(tipd_WADDR4));
   VitalWireDelay (WADDR5_ipd, WADDR5, VitalExtendToFillDelay(tipd_WADDR5));
   VitalWireDelay (WADDR6_ipd, WADDR6, VitalExtendToFillDelay(tipd_WADDR6));
   VitalWireDelay (WADDR7_ipd, WADDR7, VitalExtendToFillDelay(tipd_WADDR7));
   VitalWireDelay (RADDR0_ipd, RADDR0, VitalExtendToFillDelay(tipd_RADDR0));
   VitalWireDelay (RADDR1_ipd, RADDR1, VitalExtendToFillDelay(tipd_RADDR1));
   VitalWireDelay (RADDR2_ipd, RADDR2, VitalExtendToFillDelay(tipd_RADDR2));
   VitalWireDelay (RADDR3_ipd, RADDR3, VitalExtendToFillDelay(tipd_RADDR3));
   VitalWireDelay (RADDR4_ipd, RADDR4, VitalExtendToFillDelay(tipd_RADDR4));
   VitalWireDelay (RADDR5_ipd, RADDR5, VitalExtendToFillDelay(tipd_RADDR5));
   VitalWireDelay (RADDR6_ipd, RADDR6, VitalExtendToFillDelay(tipd_RADDR6));
   VitalWireDelay (RADDR7_ipd, RADDR7, VitalExtendToFillDelay(tipd_RADDR7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

---------------------------------------------------------------
--                  Behavior Section                         --
---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);
    WBdlyd      <= WBint after 1 ps;


    PROCESS
    BEGIN
      INIT_MEM <= '1';
      WAIT;
    END PROCESS;

    VITALBehavior : process (INIT_MEM, 
                          RADDR0_ipd, RADDR1_ipd, RADDR2_ipd, RADDR3_ipd, RADDR4_ipd, RADDR5_ipd, RADDR6_ipd, RADDR7_ipd, 
                          WADDR0_ipd, WADDR1_ipd, WADDR2_ipd, WADDR3_ipd, WADDR4_ipd, WADDR5_ipd, WADDR6_ipd, WADDR7_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd 
                          )

    -- some internal veriable declaration
     variable RAM_di_int         : std_logic_vector(8 downto 0);
     variable memory_array       : MEM_TYPE := (others =>(others => 'X'));
     variable do_par             : std_logic:= 'X';
     variable tmp_par            : std_logic:= 'X';
     variable tmp_par2           : std_logic:= 'X';
     variable wpe_var            : std_logic:= 'X';

     --  Read Timing Check Results
     variable PeriodData_RDB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RDB                  : X01                 := '0';
     variable PeriodData_RBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RBLKB                : X01                  := '0';
     variable PeriodData_RADDR0          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR0               : X01                 := '0';
     variable PeriodData_RADDR1          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR1               : X01                 := '0';
     variable PeriodData_RADDR2          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR2               : X01                 := '0';
     variable PeriodData_RADDR3          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR3               : X01                 := '0';
     variable PeriodData_RADDR4          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR4               : X01                 := '0';
     variable PeriodData_RADDR5          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR5               : X01                 := '0';
     variable PeriodData_RADDR6          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR6               : X01                 := '0';
     variable PeriodData_RADDR7          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR7               : X01                 := '0';
     variable Tviol_WADDR0_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR0_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR0_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR0_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR0_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR1_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR1_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR1_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR1_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR2_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR2_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR2_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR2_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR3_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR3_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR3_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR3_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR4_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR4_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR4_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR4_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR5_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR5_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR5_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR5_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR6_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR6_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR6_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR6_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR7_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR7_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR7_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR7_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WRB_posedge      : X01                 := '0';
     variable TmDt_DI0_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI0_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WRB_posedge      : X01                 := '0';
     variable TmDt_DI1_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI1_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WRB_posedge      : X01                 := '0';
     variable TmDt_DI2_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI2_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WRB_posedge      : X01                 := '0';
     variable TmDt_DI3_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI3_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WRB_posedge      : X01                 := '0';
     variable TmDt_DI4_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI4_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WRB_posedge      : X01                 := '0';
     variable TmDt_DI5_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI5_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WRB_posedge      : X01                 := '0';
     variable TmDt_DI6_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI6_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WRB_posedge      : X01                 := '0';
     variable TmDt_DI7_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI7_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WRB_posedge      : X01                 := '0';
     variable TmDt_DI8_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI8_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WRB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WRB                  : X01                 := '0';
     variable PeriodData_WBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WBLKB                : X01                 := '0';
     variable Tviol_RDB_WRB_posedge      : X01                 := '0';
     variable TmDt_RDB_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_WRB_negedge      : X01                 := '0';
     variable TmDt_RDB_WRB_negedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_WRB_posedge    : X01                 := '0';
     variable TmDt_RBLKB_WRB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_WRB_negedge    : X01                 := '0';
     variable TmDt_RBLKB_WRB_negedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR0_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR0_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR0_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR0_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR1_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR1_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR2_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR2_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR3_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR3_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR4_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR4_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR5_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR5_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR6_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR6_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_WRB_posedge   : X01                 := '0';
     variable TmDt_RADDR7_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_WRB_negedge   : X01                 := '0';
     variable TmDt_RADDR7_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_WBLKB_posedge    : X01                 := '0';
     variable TmDt_RDB_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_WBLKB_negedge    : X01                 := '0';
     variable TmDt_RDB_WBLKB_negedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_WBLKB_posedge  : X01                 := '0';
     variable TmDt_RBLKB_WBLKB_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_WBLKB_negedge  : X01                 := '0';
     variable TmDt_RBLKB_WBLKB_negedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR0_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR0_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR0_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR0_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR1_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR1_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR2_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR2_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR3_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR3_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR4_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR4_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR5_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR5_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR6_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR6_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_WBLKB_posedge : X01                 := '0';
     variable TmDt_RADDR7_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_WBLKB_negedge : X01                 := '0';
     variable TmDt_RADDR7_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results

     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     variable DO0_zd : std_ulogic;
     variable DO1_zd : std_ulogic;
     variable DO2_zd : std_ulogic;
     variable DO3_zd : std_ulogic;
     variable DO4_zd : std_ulogic;
     variable DO5_zd : std_ulogic;
     variable DO6_zd : std_ulogic;
     variable DO7_zd : std_ulogic;
     variable DO8_zd : std_ulogic;
     variable RPE_zd : std_ulogic;
     variable WPE_zd : std_ulogic;
     variable DOS_zd : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData  : VitalGlitchDataType;
     variable DO1_GlitchData  : VitalGlitchDataType;
     variable DO2_GlitchData  : VitalGlitchDataType;
     variable DO3_GlitchData  : VitalGlitchDataType;
     variable DO4_GlitchData  : VitalGlitchDataType;
     variable DO5_GlitchData  : VitalGlitchDataType;
     variable DO6_GlitchData  : VitalGlitchDataType;
     variable DO7_GlitchData  : VitalGlitchDataType;
     variable DO8_GlitchData  : VitalGlitchDataType;
     variable DOS_GlitchData  : VitalGlitchDataType;

     -- last value variables
     variable RBint_previous  : std_ulogic := 'X';
     variable WBint_previous  : std_ulogic := 'X';
     variable DIS_previous    : std_ulogic := 'X';
     variable RADDR0_previous : std_ulogic := 'X';
     variable RADDR1_previous : std_ulogic := 'X';
     variable RADDR2_previous : std_ulogic := 'X';
     variable RADDR3_previous : std_ulogic := 'X';
     variable RADDR4_previous : std_ulogic := 'X';
     variable RADDR5_previous : std_ulogic := 'X';
     variable RADDR6_previous : std_ulogic := 'X';
     variable RADDR7_previous : std_ulogic := 'X';
     variable WADDR0_previous : std_ulogic := 'X';
     variable WADDR1_previous : std_ulogic := 'X';
     variable WADDR2_previous : std_ulogic := 'X';
     variable WADDR3_previous : std_ulogic := 'X';
     variable WADDR4_previous : std_ulogic := 'X';
     variable WADDR5_previous : std_ulogic := 'X';
     variable WADDR6_previous : std_ulogic := 'X';
     variable WADDR7_previous : std_ulogic := 'X';

     variable PARODD_previous : std_ulogic := 'X';
     variable Write_OK        : Boolean := FALSE;

     variable inline    : LINE;
     variable indata    : std_logic_vector(8 downto 0);
     variable resdata   : std_logic_vector(8 downto 0);
     variable i         : integer:=0;
     file     memfile   : text;
     variable status         : file_open_status;

 begin -- process VITALBehavior

  -----------------------------------------------------------
  --    Initialize memory file from MEMORYFILE string      --
  -----------------------------------------------------------

  if ( INIT_MEM'EVENT and INIT_MEM = '1') then
    file_open(status, memfile, MEMORYFILE, read_mode);
    if ( status=open_ok ) then
      while((i < 256) and (not ENDFILE(memfile))) loop
        readline(memfile,inline);
        read(inline,indata);
        resdata := indata;
        memory_array(i) := resdata;
        i := i+1;
      end loop;
    else
      assert ( MEMORYFILE'length = 0 )
        report "Failed to open RAM256x9AAP memory initialization file in read mode"
        severity Note;
    end if;
    file_close(memfile);
  end if;


      WADDR := ((INT(WADDR7_ipd)*128)+(INT(WADDR6_ipd)*64)+(INT(
               WADDR5_ipd)*32) + (INT(WADDR4_ipd)*16) + 
               (INT(WADDR3_ipd)*8) + (INT(WADDR2_ipd)*4) + (INT(
               WADDR1_ipd)*2) + (INT(WADDR0_ipd)*1));
   -- Convert Read Address Signal to Integer

      RADDR := ((INT(RADDR7_ipd)*128)+(INT(RADDR6_ipd)*64)+(INT(
               RADDR5_ipd)*32) + (INT(RADDR4_ipd)*16) + 
               (INT(RADDR3_ipd)*8) + (INT(RADDR2_ipd)*4) + (INT(
               RADDR1_ipd)*2) + (INT(RADDR0_ipd)*1));

   if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

      VitalPeriodPulseCheck ( Pviol_RDB,
                              PeriodData_RDB,
                              RDB_ipd, "RDB",
                              0.0 ns,
                              tperiod_RDB,
                              tpw_RDB_posedge,
                              tpw_RDB_negedge,
                              (To_X01(RBLKB_ipd) = '0'),
                             InstancePath &"/RAM256x9AAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RBLKB,
                              PeriodData_RBLKB,
                              RBLKB_ipd, "RBLKB",
                              0.0 ns,
                              tperiod_RBLKB,
                              tpw_RBLKB_posedge,
                              tpw_RBLKB_negedge,
                              (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR0,
                              PeriodData_RADDR0,
                              RADDR0_ipd, "RADDR0",
                              0.0 ns,
                              tpw_RADDR0_posedge + tpw_RADDR0_posedge,
                              tpw_RADDR0_posedge,
                              tpw_RADDR0_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR1,
                              PeriodData_RADDR1,
                              RADDR1_ipd, "RADDR1",
                              0.0 ns,
                              tpw_RADDR1_posedge + tpw_RADDR1_posedge,
                              tpw_RADDR1_posedge,
                              tpw_RADDR1_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR2,
                              PeriodData_RADDR2,
                              RADDR2_ipd, "RADDR2",
                              0.0 ns,
                              tpw_RADDR2_posedge + tpw_RADDR2_posedge,
                              tpw_RADDR2_posedge,
                              tpw_RADDR2_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR3,
                              PeriodData_RADDR3,
                              RADDR3_ipd, "RADDR3",
                              0.0 ns,
                              tpw_RADDR3_posedge + tpw_RADDR3_posedge,
                              tpw_RADDR3_posedge,
                              tpw_RADDR3_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR4,
                              PeriodData_RADDR4,
                              RADDR4_ipd, "RADDR4",
                              0.0 ns,
                              tpw_RADDR4_posedge + tpw_RADDR4_posedge,
                              tpw_RADDR4_posedge,
                              tpw_RADDR4_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR5,
                              PeriodData_RADDR5,
                              RADDR5_ipd, "RADDR5",
                              0.0 ns,
                              tpw_RADDR5_posedge + tpw_RADDR5_posedge,
                              tpw_RADDR5_posedge,
                              tpw_RADDR5_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR6,
                              PeriodData_RADDR6,
                              RADDR6_ipd, "RADDR6",
                              0.0 ns,
                              tpw_RADDR6_posedge + tpw_RADDR6_posedge,
                              tpw_RADDR6_posedge,
                              tpw_RADDR6_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR7,
                              PeriodData_RADDR7,
                              RADDR7_ipd, "RADDR7",
                              0.0 ns,
                              tpw_RADDR7_posedge + tpw_RADDR7_posedge,
                              tpw_RADDR7_posedge,
                              tpw_RADDR7_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AAP",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_negedge,
                             TmDt_WADDR0_WRB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR0_WRB_posedge_negedge,
                             tsetup_WADDR0_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_negedge,
                             TmDt_WADDR0_WRB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR0_WRB_negedge_negedge,
                             tsetup_WADDR0_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_negedge,
                             TmDt_WADDR1_WRB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR1_WRB_posedge_negedge,
                             tsetup_WADDR1_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_negedge,
                             TmDt_WADDR1_WRB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR1_WRB_negedge_negedge,
                             tsetup_WADDR1_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_negedge,
                             TmDt_WADDR2_WRB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR2_WRB_posedge_negedge,
                             tsetup_WADDR2_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_negedge,
                             TmDt_WADDR2_WRB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR2_WRB_negedge_negedge,
                             tsetup_WADDR2_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_negedge,
                             TmDt_WADDR3_WRB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR3_WRB_posedge_negedge,
                             tsetup_WADDR3_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_negedge,
                             TmDt_WADDR3_WRB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR3_WRB_negedge_negedge,
                             tsetup_WADDR3_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_negedge,
                             TmDt_WADDR4_WRB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR4_WRB_posedge_negedge,
                             tsetup_WADDR4_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_negedge,
                             TmDt_WADDR4_WRB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR4_WRB_negedge_negedge,
                             tsetup_WADDR4_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_negedge,
                             TmDt_WADDR5_WRB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR5_WRB_posedge_negedge,
                             tsetup_WADDR5_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_negedge,
                             TmDt_WADDR5_WRB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR5_WRB_negedge_negedge,
                             tsetup_WADDR5_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_negedge,
                             TmDt_WADDR6_WRB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR6_WRB_posedge_negedge,
                             tsetup_WADDR6_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_negedge,
                             TmDt_WADDR6_WRB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR6_WRB_negedge_negedge,
                             tsetup_WADDR6_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_negedge,
                             TmDt_WADDR7_WRB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR7_WRB_posedge_negedge,
                             tsetup_WADDR7_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_negedge,
                             TmDt_WADDR7_WRB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR7_WRB_negedge_negedge,
                             tsetup_WADDR7_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_negedge,
                             TmDt_WADDR0_WBLKB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR0_WBLKB_posedge_negedge,
                             tsetup_WADDR0_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_negedge,
                             TmDt_WADDR0_WBLKB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR0_WBLKB_negedge_negedge,
                             tsetup_WADDR0_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_negedge,
                             TmDt_WADDR1_WBLKB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR1_WBLKB_posedge_negedge,
                             tsetup_WADDR1_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_negedge,
                             TmDt_WADDR1_WBLKB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR1_WBLKB_negedge_negedge,
                             tsetup_WADDR1_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_negedge,
                             TmDt_WADDR2_WBLKB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR2_WBLKB_posedge_negedge,
                             tsetup_WADDR2_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_negedge,
                             TmDt_WADDR2_WBLKB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR2_WBLKB_negedge_negedge,
                             tsetup_WADDR2_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_negedge,
                             TmDt_WADDR3_WBLKB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR3_WBLKB_posedge_negedge,
                             tsetup_WADDR3_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_negedge,
                             TmDt_WADDR3_WBLKB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR3_WBLKB_negedge_negedge,
                             tsetup_WADDR3_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_negedge,
                             TmDt_WADDR4_WBLKB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR4_WBLKB_posedge_negedge,
                             tsetup_WADDR4_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_negedge,
                             TmDt_WADDR4_WBLKB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR4_WBLKB_negedge_negedge,
                             tsetup_WADDR4_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_negedge,
                             TmDt_WADDR5_WBLKB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR5_WBLKB_posedge_negedge,
                             tsetup_WADDR5_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_negedge,
                             TmDt_WADDR5_WBLKB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR5_WBLKB_negedge_negedge,
                             tsetup_WADDR5_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_negedge,
                             TmDt_WADDR6_WBLKB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR6_WBLKB_posedge_negedge,
                             tsetup_WADDR6_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_negedge,
                             TmDt_WADDR6_WBLKB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR6_WBLKB_negedge_negedge,
                             tsetup_WADDR6_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_negedge,
                             TmDt_WADDR7_WBLKB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR7_WBLKB_posedge_negedge,
                             tsetup_WADDR7_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_negedge,
                             TmDt_WADDR7_WBLKB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR7_WBLKB_negedge_negedge,
                             tsetup_WADDR7_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_posedge,
                             TmDt_WADDR0_WRB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WRB_posedge_posedge,
                             thold_WADDR0_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_posedge,
                             TmDt_WADDR0_WRB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WRB_negedge_posedge,
                             thold_WADDR0_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_posedge,
                             TmDt_WADDR1_WRB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WRB_posedge_posedge,
                             thold_WADDR1_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_posedge,
                             TmDt_WADDR1_WRB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WRB_negedge_posedge,
                             thold_WADDR1_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_posedge,
                             TmDt_WADDR2_WRB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WRB_posedge_posedge,
                             thold_WADDR2_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_posedge,
                             TmDt_WADDR2_WRB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WRB_negedge_posedge,
                             thold_WADDR2_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_posedge,
                             TmDt_WADDR3_WRB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WRB_posedge_posedge,
                             thold_WADDR3_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_posedge,
                             TmDt_WADDR3_WRB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WRB_negedge_posedge,
                             thold_WADDR3_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_posedge,
                             TmDt_WADDR4_WRB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WRB_posedge_posedge,
                             thold_WADDR4_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_posedge,
                             TmDt_WADDR4_WRB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WRB_negedge_posedge,
                             thold_WADDR4_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_posedge,
                             TmDt_WADDR5_WRB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WRB_posedge_posedge,
                             thold_WADDR5_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_posedge,
                             TmDt_WADDR5_WRB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WRB_negedge_posedge,
                             thold_WADDR5_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_posedge,
                             TmDt_WADDR6_WRB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WRB_posedge_posedge,
                             thold_WADDR6_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_posedge,
                             TmDt_WADDR6_WRB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WRB_negedge_posedge,
                             thold_WADDR6_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_posedge,
                             TmDt_WADDR7_WRB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WRB_posedge_posedge,
                             thold_WADDR7_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_posedge,
                             TmDt_WADDR7_WRB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WRB_negedge_posedge,
                             thold_WADDR7_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_posedge,
                             TmDt_WADDR0_WBLKB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WBLKB_posedge_posedge,
                             thold_WADDR0_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_posedge,
                             TmDt_WADDR0_WBLKB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WBLKB_negedge_posedge,
                             thold_WADDR0_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_posedge,
                             TmDt_WADDR1_WBLKB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WBLKB_posedge_posedge,
                             thold_WADDR1_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_posedge,
                             TmDt_WADDR1_WBLKB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WBLKB_negedge_posedge,
                             thold_WADDR1_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_posedge,
                             TmDt_WADDR2_WBLKB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WBLKB_posedge_posedge,
                             thold_WADDR2_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_posedge,
                             TmDt_WADDR2_WBLKB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WBLKB_negedge_posedge,
                             thold_WADDR2_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_posedge,
                             TmDt_WADDR3_WBLKB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WBLKB_posedge_posedge,
                             thold_WADDR3_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_posedge,
                             TmDt_WADDR3_WBLKB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WBLKB_negedge_posedge,
                             thold_WADDR3_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_posedge,
                             TmDt_WADDR4_WBLKB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WBLKB_posedge_posedge,
                             thold_WADDR4_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_posedge,
                             TmDt_WADDR4_WBLKB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WBLKB_negedge_posedge,
                             thold_WADDR4_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_posedge,
                             TmDt_WADDR5_WBLKB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WBLKB_posedge_posedge,
                             thold_WADDR5_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_posedge,
                             TmDt_WADDR5_WBLKB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WBLKB_negedge_posedge,
                             thold_WADDR5_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_posedge,
                             TmDt_WADDR6_WBLKB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WBLKB_posedge_posedge,
                             thold_WADDR6_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_posedge,
                             TmDt_WADDR6_WBLKB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WBLKB_negedge_posedge,
                             thold_WADDR6_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_posedge,
                             TmDt_WADDR7_WBLKB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WBLKB_posedge_posedge,
                             thold_WADDR7_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_posedge,
                             TmDt_WADDR7_WBLKB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WBLKB_negedge_posedge,
                             thold_WADDR7_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_posedge_posedge,
                             tsetup_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_negedge_posedge,
                             tsetup_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_posedge_posedge,
                             tsetup_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_negedge_posedge,
                             tsetup_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_posedge_posedge,
                             tsetup_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_negedge_posedge,
                             tsetup_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_posedge_posedge,
                             tsetup_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_negedge_posedge,
                             tsetup_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_posedge_posedge,
                             tsetup_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_negedge_posedge,
                             tsetup_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_posedge_posedge,
                             tsetup_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_negedge_posedge,
                             tsetup_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_posedge_posedge,
                             tsetup_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_negedge_posedge,
                             tsetup_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_posedge_posedge,
                             tsetup_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_negedge_posedge,
                             tsetup_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_posedge_posedge,
                             tsetup_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_negedge_posedge,
                             tsetup_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_posedge_posedge,
                             tsetup_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_negedge_posedge,
                             tsetup_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_posedge_posedge,
                             tsetup_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_negedge_posedge,
                             tsetup_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_posedge_posedge,
                             tsetup_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_negedge_posedge,
                             tsetup_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_posedge_posedge,
                             tsetup_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_negedge_posedge,
                             tsetup_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_posedge_posedge,
                             tsetup_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_negedge_posedge,
                             tsetup_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_posedge_posedge,
                             tsetup_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_negedge_posedge,
                             tsetup_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_posedge_posedge,
                             tsetup_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_negedge_posedge,
                             tsetup_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_posedge_posedge,
                             tsetup_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_negedge_posedge,
                             tsetup_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_posedge_posedge,
                             tsetup_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_negedge_posedge,
                             tsetup_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AAP",
                             True,
                             True,
                             WARNING
                             );
      VitalPeriodPulseCheck ( Pviol_WBLKB,
                              PeriodData_WBLKB,
                              WBLKB_ipd, "WBLKB",
                              0.0 ns,
                              tperiod_WBLKB,
                              tpw_WBLKB_posedge,
                              tpw_WBLKB_negedge,
                              (To_X01(WRB_ipd) = '0'),
                              InstancePath & "/RAM256x9AAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_WRB,
                              PeriodData_WRB,
                              WRB_ipd, "WRB",
                              0.0 ns,
                              tperiod_WRB,
                              tpw_WRB_posedge,
                              tpw_WRB_negedge,
                              (To_X01(WBLKB_ipd) = '0'),
                              InstancePath & "/RAM256x9AAP",
                              True,
                              True,
                              WARNING
                              );
   ------------------------------------------------------------
   --        Timing Checking for Read and write conflict     --
   ------------------------------------------------------------
       VitalSetupHoldCheck ( Tviol_RDB_WRB_negedge,
                             TmDt_RDB_WRB_negedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_RDB_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_WBLKB_negedge,
                             TmDt_RDB_WBLKB_negedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_RDB_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB) = '0') AND (To_X01(RBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_WRB_posedge,
                             TmDt_RDB_WRB_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RDB_WRB_posedge_posedge,
                             0.0 ns,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_WBLKB_posedge,
                             TmDt_RDB_WBLKB_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RDB_WBLKB_posedge_posedge,
                             0.0 ns,
                             (To_X01(WRB) = '0') AND (To_X01(RBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_WRB_negedge,
                             TmDt_RBLKB_WRB_negedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_RBLKB_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB) = '0') AND (To_X01(RDB_ipd) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_WBLKB_negedge,
                             TmDt_RBLKB_WBLKB_negedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_RBLKB_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB) = '0') AND (To_X01(RDB_ipd) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_WRB_posedge,
                             TmDt_RBLKB_WRB_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RBLKB_WRB_posedge_posedge,
                             0.0 ns,
                             (To_X01(WBLKB) = '0') AND (To_X01(RDB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_WBLKB_posedge,
                             TmDt_RBLKB_WBLKB_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RBLKB_WBLKB_posedge_posedge,
                             0.0 ns,
                             (To_X01(WRB) = '0') AND (To_X01(RDB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WRB_posedge,
                             TmDt_RADDR0_WRB_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR0_WRB_negedge_posedge,
                             thold_RADDR0_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WRB_posedge,
                             TmDt_RADDR0_WRB_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR0_WRB_posedge_posedge,
                             thold_RADDR0_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WRB_negedge,
                             TmDt_RADDR0_WRB_negedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR0_WRB_posedge_negedge,
                             tsetup_RADDR0_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WRB_negedge,
                             TmDt_RADDR0_WRB_negedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR0_WRB_negedge_negedge,
                             tsetup_RADDR0_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WBLKB_posedge,
                             TmDt_RADDR0_WBLKB_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR0_WRB_negedge_posedge,
                             thold_RADDR0_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WBLKB_posedge,
                             TmDt_RADDR0_WBLKB_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR0_WRB_posedge_posedge,
                             thold_RADDR0_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WBLKB_negedge,
                             TmDt_RADDR0_WBLKB_negedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR0_WBLKB_posedge_negedge,
                             tsetup_RADDR0_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WBLKB_negedge,
                             TmDt_RADDR0_WBLKB_negedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR0_WBLKB_negedge_negedge,
                             tsetup_RADDR0_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WRB_posedge,
                             TmDt_RADDR1_WRB_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR1_WRB_negedge_posedge,
                             thold_RADDR1_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WRB_posedge,
                             TmDt_RADDR1_WRB_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR1_WRB_posedge_posedge,
                             thold_RADDR1_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WRB_negedge,
                             TmDt_RADDR1_WRB_negedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR1_WRB_posedge_negedge,
                             tsetup_RADDR1_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WRB_negedge,
                             TmDt_RADDR1_WRB_negedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR1_WRB_negedge_negedge,
                             tsetup_RADDR1_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WBLKB_posedge,
                             TmDt_RADDR1_WBLKB_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR1_WRB_negedge_posedge,
                             thold_RADDR1_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WBLKB_posedge,
                             TmDt_RADDR1_WBLKB_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR1_WRB_posedge_posedge,
                             thold_RADDR1_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WBLKB_negedge,
                             TmDt_RADDR1_WBLKB_negedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR1_WBLKB_posedge_negedge,
                             tsetup_RADDR1_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WBLKB_negedge,
                             TmDt_RADDR1_WBLKB_negedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR1_WBLKB_negedge_negedge,
                             tsetup_RADDR1_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WRB_posedge,
                             TmDt_RADDR2_WRB_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR2_WRB_negedge_posedge,
                             thold_RADDR2_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WRB_posedge,
                             TmDt_RADDR2_WRB_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR2_WRB_posedge_posedge,
                             thold_RADDR2_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WRB_negedge,
                             TmDt_RADDR2_WRB_negedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR2_WRB_posedge_negedge,
                             tsetup_RADDR2_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WRB_negedge,
                             TmDt_RADDR2_WRB_negedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR2_WRB_negedge_negedge,
                             tsetup_RADDR2_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WBLKB_posedge,
                             TmDt_RADDR2_WBLKB_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR2_WRB_negedge_posedge,
                             thold_RADDR2_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WBLKB_posedge,
                             TmDt_RADDR2_WBLKB_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR2_WRB_posedge_posedge,
                             thold_RADDR2_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WBLKB_negedge,
                             TmDt_RADDR2_WBLKB_negedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR2_WBLKB_posedge_negedge,
                             tsetup_RADDR2_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WBLKB_negedge,
                             TmDt_RADDR2_WBLKB_negedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR2_WBLKB_negedge_negedge,
                             tsetup_RADDR2_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WRB_posedge,
                             TmDt_RADDR3_WRB_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR3_WRB_negedge_posedge,
                             thold_RADDR3_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WRB_posedge,
                             TmDt_RADDR3_WRB_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR3_WRB_posedge_posedge,
                             thold_RADDR3_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WRB_negedge,
                             TmDt_RADDR3_WRB_negedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR3_WRB_posedge_negedge,
                             tsetup_RADDR3_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WRB_negedge,
                             TmDt_RADDR3_WRB_negedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR3_WRB_negedge_negedge,
                             tsetup_RADDR3_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WBLKB_posedge,
                             TmDt_RADDR3_WBLKB_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR3_WRB_negedge_posedge,
                             thold_RADDR3_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WBLKB_posedge,
                             TmDt_RADDR3_WBLKB_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR3_WRB_posedge_posedge,
                             thold_RADDR3_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WBLKB_negedge,
                             TmDt_RADDR3_WBLKB_negedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR3_WBLKB_posedge_negedge,
                             tsetup_RADDR3_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WBLKB_negedge,
                             TmDt_RADDR3_WBLKB_negedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR3_WBLKB_negedge_negedge,
                             tsetup_RADDR3_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WRB_posedge,
                             TmDt_RADDR4_WRB_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR4_WRB_negedge_posedge,
                             thold_RADDR4_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WRB_posedge,
                             TmDt_RADDR4_WRB_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR4_WRB_posedge_posedge,
                             thold_RADDR4_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WRB_negedge,
                             TmDt_RADDR4_WRB_negedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR4_WRB_posedge_negedge,
                             tsetup_RADDR4_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WRB_negedge,
                             TmDt_RADDR4_WRB_negedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR4_WRB_negedge_negedge,
                             tsetup_RADDR4_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WBLKB_posedge,
                             TmDt_RADDR4_WBLKB_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR4_WRB_negedge_posedge,
                             thold_RADDR4_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WBLKB_posedge,
                             TmDt_RADDR4_WBLKB_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR4_WRB_posedge_posedge,
                             thold_RADDR4_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WBLKB_negedge,
                             TmDt_RADDR4_WBLKB_negedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR4_WBLKB_posedge_negedge,
                             tsetup_RADDR4_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WBLKB_negedge,
                             TmDt_RADDR4_WBLKB_negedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR4_WBLKB_negedge_negedge,
                             tsetup_RADDR4_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WRB_posedge,
                             TmDt_RADDR5_WRB_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR5_WRB_negedge_posedge,
                             thold_RADDR5_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WRB_posedge,
                             TmDt_RADDR5_WRB_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR5_WRB_posedge_posedge,
                             thold_RADDR5_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WRB_negedge,
                             TmDt_RADDR5_WRB_negedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR5_WRB_posedge_negedge,
                             tsetup_RADDR5_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WRB_negedge,
                             TmDt_RADDR5_WRB_negedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR5_WRB_negedge_negedge,
                             tsetup_RADDR5_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WBLKB_posedge,
                             TmDt_RADDR5_WBLKB_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR5_WRB_negedge_posedge,
                             thold_RADDR5_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WBLKB_posedge,
                             TmDt_RADDR5_WBLKB_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR5_WRB_posedge_posedge,
                             thold_RADDR5_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WBLKB_negedge,
                             TmDt_RADDR5_WBLKB_negedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR5_WBLKB_posedge_negedge,
                             tsetup_RADDR5_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WBLKB_negedge,
                             TmDt_RADDR5_WBLKB_negedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR5_WBLKB_negedge_negedge,
                             tsetup_RADDR5_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WRB_posedge,
                             TmDt_RADDR6_WRB_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR6_WRB_negedge_posedge,
                             thold_RADDR6_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WRB_posedge,
                             TmDt_RADDR6_WRB_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR6_WRB_posedge_posedge,
                             thold_RADDR6_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WRB_negedge,
                             TmDt_RADDR6_WRB_negedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR6_WRB_posedge_negedge,
                             tsetup_RADDR6_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WRB_negedge,
                             TmDt_RADDR6_WRB_negedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR6_WRB_negedge_negedge,
                             tsetup_RADDR6_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WBLKB_posedge,
                             TmDt_RADDR6_WBLKB_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR6_WRB_negedge_posedge,
                             thold_RADDR6_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WBLKB_posedge,
                             TmDt_RADDR6_WBLKB_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR6_WRB_posedge_posedge,
                             thold_RADDR6_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WBLKB_negedge,
                             TmDt_RADDR6_WBLKB_negedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR6_WBLKB_posedge_negedge,
                             tsetup_RADDR6_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WBLKB_negedge,
                             TmDt_RADDR6_WBLKB_negedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR6_WBLKB_negedge_negedge,
                             tsetup_RADDR6_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WRB_posedge,
                             TmDt_RADDR7_WRB_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR7_WRB_negedge_posedge,
                             thold_RADDR7_WRB_negedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WRB_posedge,
                             TmDt_RADDR7_WRB_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR7_WRB_posedge_posedge,
                             thold_RADDR7_WRB_posedge_posedge,
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WRB_negedge,
                             TmDt_RADDR7_WRB_negedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR7_WRB_posedge_negedge,
                             tsetup_RADDR7_WRB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WRB_negedge,
                             TmDt_RADDR7_WRB_negedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_RADDR7_WRB_negedge_negedge,
                             tsetup_RADDR7_WRB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBLKB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WBLKB_posedge,
                             TmDt_RADDR7_WBLKB_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR7_WRB_negedge_posedge,
                             thold_RADDR7_WRB_negedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WBLKB_posedge,
                             TmDt_RADDR7_WBLKB_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR7_WRB_posedge_posedge,
                             thold_RADDR7_WRB_posedge_posedge,
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WBLKB_negedge,
                             TmDt_RADDR7_WBLKB_negedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR7_WBLKB_posedge_negedge,
                             tsetup_RADDR7_WBLKB_posedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WBLKB_negedge,
                             TmDt_RADDR7_WBLKB_negedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_RADDR7_WBLKB_negedge_negedge,
                             tsetup_RADDR7_WBLKB_negedge_negedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WRB) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                             InstancePath & "/ RAM256x9",
                             True,
                             True,
                             WARNING
                             );

   end if;

   ------------------------------------------------------------
   --         WPE generating  block                            -
   ------------------------------------------------------------

      tmp_par  := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;

      if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
          ( TO_X01 ( DI7_ipd )    = 'X' ) or
          ( TO_X01 ( DI6_ipd )    = 'X' ) or
          ( TO_X01 ( DI5_ipd )    = 'X' ) or
          ( TO_X01 ( DI4_ipd )    = 'X' ) or
          ( TO_X01 ( DI3_ipd )    = 'X' ) or
          ( TO_X01 ( DI2_ipd )    = 'X' ) or
          ( TO_X01 ( DI1_ipd )    = 'X' ) or
          ( TO_X01 ( DI0_ipd )    = 'X' )
         ) then
        wpe_var  :=  'X';
      else
        if ( tmp_par /= PARODD_ipd ) then
          wpe_var  :=  '1';
        else
          wpe_var  :=  '0';
        end if;
      end if;
      RAM_di_int(8) := wpe_var;
      WPE_zd := wpe_var;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

    if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
    end if; 

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

   if (( TO_X01 ( WBint ) = '0' ) and ( TO_X01 ( WBint_previous ) = '1' )) then
     Write_OK := True;
   end if;

 -- async memory writing 
   if ( WBint'event or WADDR0_ipd'event or WADDR1_ipd'event or 
        WADDR2_ipd'event or WADDR3_ipd'event or WADDR4_ipd'event or 
        WADDR5_ipd'event or WADDR6_ipd'event or WADDR7_ipd'event or 
        DI7_ipd'event or DI6_ipd'event or DI5_ipd'event or 
        DI4_ipd'event or DI3_ipd'event or DI2_ipd'event or 
        DI1_ipd'event or DI0_ipd'event or DI8_ipd'event ) then
     if (TO_X01(WBint)='X') then
       if (TO_X01(WBint_previous) /= 'X') then
         assert false
           report ": WRB or WBLKB unknown"
           severity Warning;
       end if;
     elsif ( TO_X01(WBint) = '0' and Write_OK ) then
          if(WADDR < 0) then
           if((TO_X01(WADDR0_ipd) = 'X') and (TO_X01(WADDR0_previous) /= 'X')) then
             assert false
             report ": WADDR0 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR1_ipd) = 'X') and (TO_X01(WADDR1_previous) /= 'X')) then
             assert false
             report ": WADDR1 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR2_ipd) = 'X') and (TO_X01(WADDR2_previous) /= 'X')) then
             assert false
             report ": WADDR2 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR3_ipd) = 'X') and (TO_X01(WADDR3_previous) /= 'X')) then
             assert false
             report ": WADDR3 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR4_ipd) = 'X') and (TO_X01(WADDR4_previous) /= 'X')) then
             assert false
             report ": WADDR4 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR5_ipd) = 'X') and (TO_X01(WADDR5_previous) /= 'X')) then
             assert false
             report ": WADDR5 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR6_ipd) = 'X') and (TO_X01(WADDR6_previous) /= 'X')) then
             assert false
             report ": WADDR6 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR7_ipd) = 'X') and (TO_X01(WADDR7_previous) /= 'X')) then
             assert false
             report ": WADDR7 unknown, no data written ......"
             severity Warning;
           end if;
          else
            RAM_di_int ( 7 downto 0 ) := DI7_ipd & DI6_ipd & DI5_ipd & DI4_ipd & 
                                          DI3_ipd & DI2_ipd & DI1_ipd & DI0_ipd;
            memory_array ( WADDR ) := RAM_di_int;
          end if;
        end if;
      end if;


 -----------------------------------------------------------
 --  Read Functional Section                              --
 -----------------------------------------------------------



-- Asynchronous RAM Read, Enable signal controlled;

   if ( RBint'event or RADDR0_ipd'event or RADDR1_ipd'event or 
        RADDR2_ipd'event or RADDR3_ipd'event or RADDR4_ipd'event or 
        RADDR5_ipd'event or RADDR6_ipd'event or RADDR7_ipd'event or
        WBint'event or WADDR0_ipd'event or WADDR1_ipd'event or 
        WADDR2_ipd'event or WADDR3_ipd'event or WADDR4_ipd'event or 
        WADDR5_ipd'event or WADDR6_ipd'event or WADDR7_ipd'event
      ) then
     if ( TO_X01 ( RBint ) = 'X' ) then
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          RPE_zd :='X';
          if (TO_X01(RBint_previous) /= 'X') then
             assert false
               report ": RDB or RBLKB unknown"
               severity Warning;
          end if;
     elsif ( RADDR < 0 ) then
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          RPE_zd :='X';
          if(TO_X01(RADDR0_ipd) = 'X') and (TO_X01(RADDR0_previous) /= 'X') then
             assert false
             report ": RADDR0 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR1_ipd) = 'X') and (TO_X01(RADDR1_previous) /= 'X') then
             assert false
             report ": RADDR1 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR2_ipd) = 'X') and (TO_X01(RADDR2_previous) /= 'X') then
             assert false
             report ": RADDR2 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR3_ipd) = 'X') and (TO_X01(RADDR3_previous) /= 'X') then
             assert false
             report ": RADDR3 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR4_ipd) = 'X') and (TO_X01(RADDR4_previous) /= 'X') then
             assert false
             report ": RADDR4 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR5_ipd) = 'X') and (TO_X01(RADDR5_previous) /= 'X') then
             assert false
             report ": RADDR5 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR6_ipd) = 'X') and (TO_X01(RADDR6_previous) /= 'X') then
             assert false
             report ": RADDR6 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR7_ipd) = 'X') and (TO_X01(RADDR7_previous) /= 'X') then
             assert false
             report ": RADDR7 unknown"
             severity Warning;
          end if;
     elsif ( WADDR = RADDR ) then
       if (( RBint'event AND ( TO_X01 ( RBint ) = '0' ) AND ( TO_X01 ( WBint ) = '1' )) OR
           ( WBint'event AND ( TO_X01 ( WBint ) = '1' ) AND ( TO_X01 ( RBint ) = '0' )) OR
           ( RBint'event AND ( TO_X01 ( RBint ) = '1' ) AND ( TO_X01 ( WBdlyd ) = '0' )) OR
           (( TO_X01 ( WBint ) = '1' ) AND ( TO_X01 ( RBint ) = '0' ) AND 
            ( RADDR0_ipd'event or RADDR1_ipd'event or 
              RADDR2_ipd'event or RADDR3_ipd'event or RADDR4_ipd'event or 
              RADDR5_ipd'event or RADDR6_ipd'event or RADDR7_ipd'event ))
          ) then
             DO0_zd := memory_array(RADDR)(0);
             DO1_zd := memory_array(RADDR)(1);
             DO2_zd := memory_array(RADDR)(2);
             DO3_zd := memory_array(RADDR)(3);
             DO4_zd := memory_array(RADDR)(4);
             DO5_zd := memory_array(RADDR)(5);
             DO6_zd := memory_array(RADDR)(6);
             DO7_zd := memory_array(RADDR)(7);
             DO8_zd := memory_array(RADDR)(8);
       end if;
     else -- WADDR /= RADDR
       if ((( TO_X01 ( WBint ) = '0' ) AND ( TO_X01 ( RBint ) = '0' ) AND
            ( RADDR0_ipd'event or RADDR1_ipd'event or RADDR2_ipd'event or 
              RADDR3_ipd'event or RADDR4_ipd'event or RADDR5_ipd'event or 
              RADDR6_ipd'event or RADDR7_ipd'event or WADDR0_ipd'event or 
              WADDR1_ipd'event or WADDR2_ipd'event or WADDR3_ipd'event or 
              WADDR4_ipd'event or WADDR5_ipd'event or WADDR6_ipd'event or 
              WADDR7_ipd'event)) OR
           ( RBint'event AND ( TO_X01 ( RBint ) = '0' )) OR
           (( TO_X01 ( RBint ) = '0' ) AND
            ( RADDR0_ipd'event or RADDR1_ipd'event or RADDR2_ipd'event or 
              RADDR3_ipd'event or RADDR4_ipd'event or RADDR5_ipd'event or 
              RADDR6_ipd'event or RADDR7_ipd'event or WADDR0_ipd'event or 
              WADDR1_ipd'event or WADDR2_ipd'event or WADDR3_ipd'event or 
              WADDR4_ipd'event or WADDR5_ipd'event or WADDR6_ipd'event or 
              WADDR7_ipd'event))
          ) then
             DO0_zd := memory_array(RADDR)(0);
             DO1_zd := memory_array(RADDR)(1);
             DO2_zd := memory_array(RADDR)(2);
             DO3_zd := memory_array(RADDR)(3);
             DO4_zd := memory_array(RADDR)(4);
             DO5_zd := memory_array(RADDR)(5);
             DO6_zd := memory_array(RADDR)(6);
             DO7_zd := memory_array(RADDR)(7);
             DO8_zd := memory_array(RADDR)(8);
       end if;
     end if;
   end if;


  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       RBint_previous  := RBint;
       WBint_previous  := WBint;
       RADDR0_previous := RADDR0_ipd;
       RADDR1_previous := RADDR1_ipd;
       RADDR2_previous := RADDR2_ipd;
       RADDR3_previous := RADDR3_ipd;
       RADDR4_previous := RADDR4_ipd;
       RADDR5_previous := RADDR5_ipd;
       RADDR6_previous := RADDR6_ipd;
       RADDR7_previous := RADDR7_ipd;
       WADDR0_previous := WADDR0_ipd;
       WADDR1_previous := WADDR1_ipd;
       WADDR2_previous := WADDR2_ipd;
       WADDR3_previous := WADDR3_ipd;
       WADDR4_previous := WADDR4_ipd;
       WADDR5_previous := WADDR5_ipd;
       WADDR6_previous := WADDR6_ipd;
       WADDR7_previous := WADDR7_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
           OutSignal     => DOS,
           GlitchData    => DOS_GlitchData,
           OutSignalName => "DOS",
           OutTemp       => DOS_zd,
           Paths  =>  (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),
           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO0), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO0), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO0), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO0), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO0), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO0), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO0), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO0), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO0), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO1), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO1), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO1), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO1), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO1), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO1), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO1), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO1), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO1), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO2), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO2), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO2), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO2), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO2), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO2), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO2), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO2), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO2), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO3), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO3), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO3), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO3), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO3), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO3), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO3), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO3), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO3), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO4), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO4), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO4), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO4), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO4), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO4), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO4), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO4), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO4), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO5), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO5), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO5), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO5), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO5), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO5), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO5), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO5), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO5), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO6), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO6), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO6), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO6), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO6), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO6), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO6), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO6), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO6), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO7), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO7), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO7), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO7), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO7), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO7), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO7), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO7), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO7), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO8), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO8), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO8), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO8), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO8), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO8), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO8), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO8), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO8), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

   end process VITALBehavior;

 end VITAL_ACT;
 
 configuration CFG_RAM256x9AA_VITAL of RAM256x9AA is
    for VITAL_ACT
    end for;
 end CFG_RAM256x9AA_VITAL;
 
 
LIBRARY ieee;
LIBRARY STD;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

USE std.textio.all;
USE ieee.std_logic_textio.all;
LIBRARY a500k;
USE a500k.all;

entity RAM256x9AST is 

   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI0_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI1_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI2_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI3_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI4_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI5_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI6_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI7_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI8_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                           : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                         : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                         : VitalDelayType := 0.000 ns;
 	tperiod_WRB                             : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WRB_RCLKS_negedge_posedge        : VitalDelayType := 0.000 ns;
 	thold_WRB_RCLKS_negedge_posedge         : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RCLKS_negedge_posedge      : VitalDelayType := 0.000 ns;
	thold_WBLKB_RCLKS_negedge_posedge       : VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';
   WPE    :  OUT STD_LOGIC := 'X';
   RPE    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');

ATTRIBUTE VITAL_LEVEL0 OF RAM256x9AST : entity IS True ;
END RAM256x9AST;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of RAM256x9AST is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal WADDR0_ipd : std_ulogic := 'X';
   signal WADDR1_ipd : std_ulogic := 'X';
   signal WADDR2_ipd : std_ulogic := 'X';
   signal WADDR3_ipd : std_ulogic := 'X';
   signal WADDR4_ipd : std_ulogic := 'X';
   signal WADDR5_ipd : std_ulogic := 'X';
   signal WADDR6_ipd : std_ulogic := 'X';
   signal WADDR7_ipd : std_ulogic := 'X';
   signal RADDR0_ipd : std_ulogic := 'X';
   signal RADDR1_ipd : std_ulogic := 'X';
   signal RADDR2_ipd : std_ulogic := 'X';
   signal RADDR3_ipd : std_ulogic := 'X';
   signal RADDR4_ipd : std_ulogic := 'X';
   signal RADDR5_ipd : std_ulogic := 'X';
   signal RADDR6_ipd : std_ulogic := 'X';
   signal RADDR7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

	-- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';
   signal INIT_MEM   : std_logic:= '0';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic:= 'X';
   signal par_f2     : std_logic:= 'X';

 begin  --  VITAL_ACT
   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (WADDR0_ipd, WADDR0, VitalExtendToFillDelay(tipd_WADDR0));
   VitalWireDelay (WADDR1_ipd, WADDR1, VitalExtendToFillDelay(tipd_WADDR1));
   VitalWireDelay (WADDR2_ipd, WADDR2, VitalExtendToFillDelay(tipd_WADDR2));
   VitalWireDelay (WADDR3_ipd, WADDR3, VitalExtendToFillDelay(tipd_WADDR3));
   VitalWireDelay (WADDR4_ipd, WADDR4, VitalExtendToFillDelay(tipd_WADDR4));
   VitalWireDelay (WADDR5_ipd, WADDR5, VitalExtendToFillDelay(tipd_WADDR5));
   VitalWireDelay (WADDR6_ipd, WADDR6, VitalExtendToFillDelay(tipd_WADDR6));
   VitalWireDelay (WADDR7_ipd, WADDR7, VitalExtendToFillDelay(tipd_WADDR7));
   VitalWireDelay (RADDR0_ipd, RADDR0, VitalExtendToFillDelay(tipd_RADDR0));
   VitalWireDelay (RADDR1_ipd, RADDR1, VitalExtendToFillDelay(tipd_RADDR1));
   VitalWireDelay (RADDR2_ipd, RADDR2, VitalExtendToFillDelay(tipd_RADDR2));
   VitalWireDelay (RADDR3_ipd, RADDR3, VitalExtendToFillDelay(tipd_RADDR3));
   VitalWireDelay (RADDR4_ipd, RADDR4, VitalExtendToFillDelay(tipd_RADDR4));
   VitalWireDelay (RADDR5_ipd, RADDR5, VitalExtendToFillDelay(tipd_RADDR5));
   VitalWireDelay (RADDR6_ipd, RADDR6, VitalExtendToFillDelay(tipd_RADDR6));
   VitalWireDelay (RADDR7_ipd, RADDR7, VitalExtendToFillDelay(tipd_RADDR7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

---------------------------------------------------------------
--                  Behavior Section                         --
---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);


    PROCESS
    BEGIN
      INIT_MEM <= '1';
      WAIT;
    END PROCESS;

    VITALBehavior : process (INIT_MEM, 
                          RADDR0_ipd, RADDR1_ipd, RADDR2_ipd, RADDR3_ipd, RADDR4_ipd, RADDR5_ipd, RADDR6_ipd, RADDR7_ipd, 
                          WADDR0_ipd, WADDR1_ipd, WADDR2_ipd, WADDR3_ipd, WADDR4_ipd, WADDR5_ipd, WADDR6_ipd, WADDR7_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd 
                          )

    -- some internal veriable declaration
     variable RAM_di_int         : std_logic_vector(8 downto 0);
     variable memory_array       : MEM_TYPE := (others =>(others => 'X'));
     variable do_par             : std_logic:= 'X';
     variable tmp_par            : std_logic:= 'X';
     variable tmp_par2           : std_logic:= 'X';
     variable wpe_var            : std_logic:= 'X';

     --  Read Timing Check Results
     variable Tviol_RADDR0_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR0_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR1_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR2_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR3_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR4_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR5_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR6_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR7_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable Tviol_WADDR0_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR0_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR0_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR0_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR0_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR1_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR1_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR1_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR1_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR2_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR2_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR2_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR2_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR3_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR3_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR3_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR3_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR4_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR4_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR4_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR4_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR5_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR5_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR5_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR5_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR6_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR6_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR6_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR6_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR7_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR7_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR7_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR7_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WRB_posedge      : X01                 := '0';
     variable TmDt_DI0_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI0_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WRB_posedge      : X01                 := '0';
     variable TmDt_DI1_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI1_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WRB_posedge      : X01                 := '0';
     variable TmDt_DI2_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI2_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WRB_posedge      : X01                 := '0';
     variable TmDt_DI3_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI3_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WRB_posedge      : X01                 := '0';
     variable TmDt_DI4_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI4_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WRB_posedge      : X01                 := '0';
     variable TmDt_DI5_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI5_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WRB_posedge      : X01                 := '0';
     variable TmDt_DI6_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI6_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WRB_posedge      : X01                 := '0';
     variable TmDt_DI7_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI7_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WRB_posedge      : X01                 := '0';
     variable TmDt_DI8_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI8_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WRB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WRB                  : X01                 := '0';
     variable PeriodData_WBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WBLKB                : X01                 := '0';
     variable Tviol_WRB_RCLKS_posedge    : X01 := '0';
     variable TmDt_WRB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_RCLKS_posedge  : X01 := '0';
     variable TmDt_WBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results

     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     variable DO0_zd : std_ulogic;
     variable DO1_zd : std_ulogic;
     variable DO2_zd : std_ulogic;
     variable DO3_zd : std_ulogic;
     variable DO4_zd : std_ulogic;
     variable DO5_zd : std_ulogic;
     variable DO6_zd : std_ulogic;
     variable DO7_zd : std_ulogic;
     variable DO8_zd : std_ulogic;
     variable RPE_zd : std_ulogic;
     variable WPE_zd : std_ulogic;
     variable DOS_zd : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData  : VitalGlitchDataType;
     variable DO1_GlitchData  : VitalGlitchDataType;
     variable DO2_GlitchData  : VitalGlitchDataType;
     variable DO3_GlitchData  : VitalGlitchDataType;
     variable DO4_GlitchData  : VitalGlitchDataType;
     variable DO5_GlitchData  : VitalGlitchDataType;
     variable DO6_GlitchData  : VitalGlitchDataType;
     variable DO7_GlitchData  : VitalGlitchDataType;
     variable DO8_GlitchData  : VitalGlitchDataType;
     variable RPE_GlitchData  : VitalGlitchDataType;
     variable WPE_GlitchData  : VitalGlitchDataType;
     variable DOS_GlitchData  : VitalGlitchDataType;

     -- last value variables
     variable RCLKS_previous  : std_ulogic := 'X';
     variable RBint_delayed   : std_ulogic := 'X';
     variable RBint_previous  : std_ulogic := 'X';
     variable WBint_previous  : std_ulogic := 'X';
     variable DIS_previous    : std_ulogic := 'X';
     variable RADDR0_delayed  : std_ulogic := 'X';
     variable RADDR1_delayed  : std_ulogic := 'X';
     variable RADDR2_delayed  : std_ulogic := 'X';
     variable RADDR3_delayed  : std_ulogic := 'X';
     variable RADDR4_delayed  : std_ulogic := 'X';
     variable RADDR5_delayed  : std_ulogic := 'X';
     variable RADDR6_delayed  : std_ulogic := 'X';
     variable RADDR7_delayed  : std_ulogic := 'X';
     variable RADDR0_previous : std_ulogic := 'X';
     variable RADDR1_previous : std_ulogic := 'X';
     variable RADDR2_previous : std_ulogic := 'X';
     variable RADDR3_previous : std_ulogic := 'X';
     variable RADDR4_previous : std_ulogic := 'X';
     variable RADDR5_previous : std_ulogic := 'X';
     variable RADDR6_previous : std_ulogic := 'X';
     variable RADDR7_previous : std_ulogic := 'X';
     variable WADDR0_previous : std_ulogic := 'X';
     variable WADDR1_previous : std_ulogic := 'X';
     variable WADDR2_previous : std_ulogic := 'X';
     variable WADDR3_previous : std_ulogic := 'X';
     variable WADDR4_previous : std_ulogic := 'X';
     variable WADDR5_previous : std_ulogic := 'X';
     variable WADDR6_previous : std_ulogic := 'X';
     variable WADDR7_previous : std_ulogic := 'X';

     variable PARODD_delayed  : std_ulogic := 'X';
     variable PARODD_previous : std_ulogic := 'X';
     variable Write_OK        : Boolean := FALSE;

     variable inline    : LINE;
     variable indata    : std_logic_vector(8 downto 0);
     variable resdata   : std_logic_vector(8 downto 0);
     variable i         : integer:=0;
     file     memfile   : text;
     variable status         : file_open_status;

 begin -- process VITALBehavior

  -----------------------------------------------------------
  --    Initialize memory file from MEMORYFILE string      --
  -----------------------------------------------------------

  if ( INIT_MEM'EVENT and INIT_MEM = '1') then
    file_open(status, memfile, MEMORYFILE, read_mode);
    if ( status=open_ok ) then
      while((i < 256) and (not ENDFILE(memfile))) loop
        readline(memfile,inline);
        read(inline,indata);
        resdata := indata;
        memory_array(i) := resdata;
        i := i+1;
      end loop;
    else
      assert ( MEMORYFILE'length = 0 )
        report "Failed to open RAM256x9AST memory initialization file in read mode"
        severity Note;
    end if;
    file_close(memfile);
  end if;


      WADDR := ((INT(WADDR7_ipd)*128)+(INT(WADDR6_ipd)*64)+(INT(
               WADDR5_ipd)*32) + (INT(WADDR4_ipd)*16) + 
               (INT(WADDR3_ipd)*8) + (INT(WADDR2_ipd)*4) + (INT(
               WADDR1_ipd)*2) + (INT(WADDR0_ipd)*1));
   -- Convert Read Address Signal to Integer
     if (RCLKS_ipd'EVENT AND RCLKS_ipd = '1') then
      RADDR := ((INT(RADDR7_delayed)*128)+(INT(RADDR6_delayed)*64)+(INT(
               RADDR5_delayed)*32) + (INT(RADDR4_delayed)*16) + 
               (INT(RADDR3_delayed)*8) + (INT(RADDR2_delayed)*4) + (INT(
               RADDR1_delayed)*2) + (INT(RADDR0_delayed)*1));
     end if;

if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

 -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9AST",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_negedge,
                             TmDt_WADDR0_WRB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR0_WRB_posedge_negedge,
                             tsetup_WADDR0_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_negedge,
                             TmDt_WADDR0_WRB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR0_WRB_negedge_negedge,
                             tsetup_WADDR0_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_negedge,
                             TmDt_WADDR1_WRB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR1_WRB_posedge_negedge,
                             tsetup_WADDR1_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_negedge,
                             TmDt_WADDR1_WRB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR1_WRB_negedge_negedge,
                             tsetup_WADDR1_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_negedge,
                             TmDt_WADDR2_WRB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR2_WRB_posedge_negedge,
                             tsetup_WADDR2_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_negedge,
                             TmDt_WADDR2_WRB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR2_WRB_negedge_negedge,
                             tsetup_WADDR2_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_negedge,
                             TmDt_WADDR3_WRB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR3_WRB_posedge_negedge,
                             tsetup_WADDR3_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_negedge,
                             TmDt_WADDR3_WRB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR3_WRB_negedge_negedge,
                             tsetup_WADDR3_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_negedge,
                             TmDt_WADDR4_WRB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR4_WRB_posedge_negedge,
                             tsetup_WADDR4_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_negedge,
                             TmDt_WADDR4_WRB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR4_WRB_negedge_negedge,
                             tsetup_WADDR4_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_negedge,
                             TmDt_WADDR5_WRB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR5_WRB_posedge_negedge,
                             tsetup_WADDR5_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_negedge,
                             TmDt_WADDR5_WRB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR5_WRB_negedge_negedge,
                             tsetup_WADDR5_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_negedge,
                             TmDt_WADDR6_WRB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR6_WRB_posedge_negedge,
                             tsetup_WADDR6_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_negedge,
                             TmDt_WADDR6_WRB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR6_WRB_negedge_negedge,
                             tsetup_WADDR6_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_negedge,
                             TmDt_WADDR7_WRB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR7_WRB_posedge_negedge,
                             tsetup_WADDR7_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_negedge,
                             TmDt_WADDR7_WRB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR7_WRB_negedge_negedge,
                             tsetup_WADDR7_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_negedge,
                             TmDt_WADDR0_WBLKB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR0_WBLKB_posedge_negedge,
                             tsetup_WADDR0_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_negedge,
                             TmDt_WADDR0_WBLKB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR0_WBLKB_negedge_negedge,
                             tsetup_WADDR0_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_negedge,
                             TmDt_WADDR1_WBLKB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR1_WBLKB_posedge_negedge,
                             tsetup_WADDR1_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_negedge,
                             TmDt_WADDR1_WBLKB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR1_WBLKB_negedge_negedge,
                             tsetup_WADDR1_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_negedge,
                             TmDt_WADDR2_WBLKB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR2_WBLKB_posedge_negedge,
                             tsetup_WADDR2_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_negedge,
                             TmDt_WADDR2_WBLKB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR2_WBLKB_negedge_negedge,
                             tsetup_WADDR2_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_negedge,
                             TmDt_WADDR3_WBLKB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR3_WBLKB_posedge_negedge,
                             tsetup_WADDR3_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_negedge,
                             TmDt_WADDR3_WBLKB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR3_WBLKB_negedge_negedge,
                             tsetup_WADDR3_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_negedge,
                             TmDt_WADDR4_WBLKB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR4_WBLKB_posedge_negedge,
                             tsetup_WADDR4_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_negedge,
                             TmDt_WADDR4_WBLKB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR4_WBLKB_negedge_negedge,
                             tsetup_WADDR4_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_negedge,
                             TmDt_WADDR5_WBLKB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR5_WBLKB_posedge_negedge,
                             tsetup_WADDR5_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_negedge,
                             TmDt_WADDR5_WBLKB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR5_WBLKB_negedge_negedge,
                             tsetup_WADDR5_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_negedge,
                             TmDt_WADDR6_WBLKB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR6_WBLKB_posedge_negedge,
                             tsetup_WADDR6_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_negedge,
                             TmDt_WADDR6_WBLKB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR6_WBLKB_negedge_negedge,
                             tsetup_WADDR6_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_negedge,
                             TmDt_WADDR7_WBLKB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR7_WBLKB_posedge_negedge,
                             tsetup_WADDR7_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_negedge,
                             TmDt_WADDR7_WBLKB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR7_WBLKB_negedge_negedge,
                             tsetup_WADDR7_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_posedge,
                             TmDt_WADDR0_WRB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WRB_posedge_posedge,
                             thold_WADDR0_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_posedge,
                             TmDt_WADDR0_WRB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WRB_negedge_posedge,
                             thold_WADDR0_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_posedge,
                             TmDt_WADDR1_WRB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WRB_posedge_posedge,
                             thold_WADDR1_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_posedge,
                             TmDt_WADDR1_WRB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WRB_negedge_posedge,
                             thold_WADDR1_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_posedge,
                             TmDt_WADDR2_WRB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WRB_posedge_posedge,
                             thold_WADDR2_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_posedge,
                             TmDt_WADDR2_WRB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WRB_negedge_posedge,
                             thold_WADDR2_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_posedge,
                             TmDt_WADDR3_WRB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WRB_posedge_posedge,
                             thold_WADDR3_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_posedge,
                             TmDt_WADDR3_WRB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WRB_negedge_posedge,
                             thold_WADDR3_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_posedge,
                             TmDt_WADDR4_WRB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WRB_posedge_posedge,
                             thold_WADDR4_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_posedge,
                             TmDt_WADDR4_WRB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WRB_negedge_posedge,
                             thold_WADDR4_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_posedge,
                             TmDt_WADDR5_WRB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WRB_posedge_posedge,
                             thold_WADDR5_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_posedge,
                             TmDt_WADDR5_WRB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WRB_negedge_posedge,
                             thold_WADDR5_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_posedge,
                             TmDt_WADDR6_WRB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WRB_posedge_posedge,
                             thold_WADDR6_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_posedge,
                             TmDt_WADDR6_WRB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WRB_negedge_posedge,
                             thold_WADDR6_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_posedge,
                             TmDt_WADDR7_WRB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WRB_posedge_posedge,
                             thold_WADDR7_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_posedge,
                             TmDt_WADDR7_WRB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WRB_negedge_posedge,
                             thold_WADDR7_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_posedge,
                             TmDt_WADDR0_WBLKB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WBLKB_posedge_posedge,
                             thold_WADDR0_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_posedge,
                             TmDt_WADDR0_WBLKB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WBLKB_negedge_posedge,
                             thold_WADDR0_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_posedge,
                             TmDt_WADDR1_WBLKB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WBLKB_posedge_posedge,
                             thold_WADDR1_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_posedge,
                             TmDt_WADDR1_WBLKB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WBLKB_negedge_posedge,
                             thold_WADDR1_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_posedge,
                             TmDt_WADDR2_WBLKB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WBLKB_posedge_posedge,
                             thold_WADDR2_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_posedge,
                             TmDt_WADDR2_WBLKB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WBLKB_negedge_posedge,
                             thold_WADDR2_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_posedge,
                             TmDt_WADDR3_WBLKB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WBLKB_posedge_posedge,
                             thold_WADDR3_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_posedge,
                             TmDt_WADDR3_WBLKB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WBLKB_negedge_posedge,
                             thold_WADDR3_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_posedge,
                             TmDt_WADDR4_WBLKB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WBLKB_posedge_posedge,
                             thold_WADDR4_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_posedge,
                             TmDt_WADDR4_WBLKB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WBLKB_negedge_posedge,
                             thold_WADDR4_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_posedge,
                             TmDt_WADDR5_WBLKB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WBLKB_posedge_posedge,
                             thold_WADDR5_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_posedge,
                             TmDt_WADDR5_WBLKB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WBLKB_negedge_posedge,
                             thold_WADDR5_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_posedge,
                             TmDt_WADDR6_WBLKB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WBLKB_posedge_posedge,
                             thold_WADDR6_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_posedge,
                             TmDt_WADDR6_WBLKB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WBLKB_negedge_posedge,
                             thold_WADDR6_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_posedge,
                             TmDt_WADDR7_WBLKB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WBLKB_posedge_posedge,
                             thold_WADDR7_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_posedge,
                             TmDt_WADDR7_WBLKB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WBLKB_negedge_posedge,
                             thold_WADDR7_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_posedge_posedge,
                             tsetup_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_negedge_posedge,
                             tsetup_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_posedge_posedge,
                             tsetup_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_negedge_posedge,
                             tsetup_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_posedge_posedge,
                             tsetup_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_negedge_posedge,
                             tsetup_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_posedge_posedge,
                             tsetup_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_negedge_posedge,
                             tsetup_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_posedge_posedge,
                             tsetup_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_negedge_posedge,
                             tsetup_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_posedge_posedge,
                             tsetup_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_negedge_posedge,
                             tsetup_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_posedge_posedge,
                             tsetup_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_negedge_posedge,
                             tsetup_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_posedge_posedge,
                             tsetup_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_negedge_posedge,
                             tsetup_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_posedge_posedge,
                             tsetup_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_negedge_posedge,
                             tsetup_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_posedge_posedge,
                             tsetup_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_negedge_posedge,
                             tsetup_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_posedge_posedge,
                             tsetup_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_negedge_posedge,
                             tsetup_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_posedge_posedge,
                             tsetup_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_negedge_posedge,
                             tsetup_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_posedge_posedge,
                             tsetup_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_negedge_posedge,
                             tsetup_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_posedge_posedge,
                             tsetup_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_negedge_posedge,
                             tsetup_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_posedge_posedge,
                             tsetup_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_negedge_posedge,
                             tsetup_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_posedge_posedge,
                             tsetup_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_negedge_posedge,
                             tsetup_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_posedge_posedge,
                             tsetup_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_negedge_posedge,
                             tsetup_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_posedge_posedge,
                             tsetup_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_negedge_posedge,
                             tsetup_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );
      VitalPeriodPulseCheck ( Pviol_WBLKB,
                              PeriodData_WBLKB,
                              WBLKB_ipd, "WBLKB",
                              0.0 ns,
                              tperiod_WBLKB,
                              tpw_WBLKB_posedge,
                              tpw_WBLKB_negedge,
                              (To_X01(WRB_ipd) = '0'),
                              InstancePath & "/RAM256x9AST",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_WRB,
                              PeriodData_WRB,
                              WRB_ipd, "WRB",
                              0.0 ns,
                              tperiod_WRB,
                              tpw_WRB_posedge,
                              tpw_WRB_negedge,
                              (To_X01(WBLKB_ipd) = '0'),
                              InstancePath & "/RAM256x9AST",
                              True,
                              True,
                              WARNING
                              );
   ------------------------------------------------------------
   --        Timing Checking for Read and write conflict     --
   ------------------------------------------------------------
       VitalSetupHoldCheck ( Tviol_WRB_RCLKS_posedge,
                             TmDt_WRB_RCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_WRB_RCLKS_negedge_posedge,
                             0.0 ns,
                             thold_WRB_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0') AND (To_X01(WBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_RCLKS_posedge,
                             TmDt_WBLKB_RCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_WBLKB_RCLKS_negedge_posedge,
                             0.0 ns,
                             thold_WBLKB_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0') AND (To_X01(WRB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9AST",
                             True,
                             True,
                             WARNING
                             );

 end if;

   ------------------------------------------------------------
   --    wpe output                                           -
   ------------------------------------------------------------

   if ( PARODD_ipd'EVENT ) then
     RPE_zd := not RPE_zd;
     WPE_zd := not WPE_zd;
   end if;

   ------------------------------------------------------------
   --         WPE checking  block                            -
   ------------------------------------------------------------

     tmp_par  := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;
     tmp_par2 := (tmp_par xor DI8_ipd);

      if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
          ( TO_X01 ( DI8_ipd )    = 'X' ) or
          ( TO_X01 ( DI7_ipd )    = 'X' ) or
          ( TO_X01 ( DI6_ipd )    = 'X' ) or
          ( TO_X01 ( DI5_ipd )    = 'X' ) or
          ( TO_X01 ( DI4_ipd )    = 'X' ) or
          ( TO_X01 ( DI3_ipd )    = 'X' ) or
          ( TO_X01 ( DI2_ipd )    = 'X' ) or
          ( TO_X01 ( DI1_ipd )    = 'X' ) or
          ( TO_X01 ( DI0_ipd )    = 'X' )
         ) then
        wpe_var  :=  'X';
      else
        if ( tmp_par2 /= PARODD_ipd ) then
          wpe_var  :=  '1';
        else
          wpe_var  :=  '0';
        end if;
      end if;
      RAM_di_int(8) := DI8_ipd;
      WPE_zd := wpe_var;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

    if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
    end if; 

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

   if (( TO_X01 ( WBint ) = '0' ) and ( TO_X01 ( WBint_previous ) = '1' )) then
     Write_OK := True;
   end if;


 -- async memory writing 
    if (TO_X01(WBint)='X') then
      if (TO_X01(WBint_previous) /= 'X') then
        assert false
        report ": WRB or WBLKB unknown"
        severity Warning;
      end if;
     elsif ( TO_X01(WBint) = '0' and Write_OK ) then
          if(WADDR < 0) then
           if((TO_X01(WADDR0_ipd) = 'X') and (TO_X01(WADDR0_previous) /= 'X')) then
             assert false
             report ": WADDR0 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR1_ipd) = 'X') and (TO_X01(WADDR1_previous) /= 'X')) then
             assert false
             report ": WADDR1 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR2_ipd) = 'X') and (TO_X01(WADDR2_previous) /= 'X')) then
             assert false
             report ": WADDR2 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR3_ipd) = 'X') and (TO_X01(WADDR3_previous) /= 'X')) then
             assert false
             report ": WADDR3 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR4_ipd) = 'X') and (TO_X01(WADDR4_previous) /= 'X')) then
             assert false
             report ": WADDR4 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR5_ipd) = 'X') and (TO_X01(WADDR5_previous) /= 'X')) then
             assert false
             report ": WADDR5 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR6_ipd) = 'X') and (TO_X01(WADDR6_previous) /= 'X')) then
             assert false
             report ": WADDR6 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR7_ipd) = 'X') and (TO_X01(WADDR7_previous) /= 'X')) then
             assert false
             report ": WADDR7 unknown, no data written ......"
             severity Warning;
           end if;
          else
             RAM_di_int(7 downto 0) :=DI7_ipd & DI6_ipd & DI5_ipd & DI4_ipd & DI3_ipd & DI2_ipd & DI1_ipd & DI0_ipd;
             memory_array(WADDR)  := RAM_di_int;
          end if;

    end if;


 -----------------------------------------------------------
 --  Read Functional Section                              --
 -----------------------------------------------------------


    if (TO_X01(RCLKS_ipd) = 'X') then
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          RPE_zd := 'X';
       if (TO_X01(RCLKS_previous) /= 'X') then
         assert false
         report ": RCLK unknown"
         severity Warning;
       end if;
    elsif(RCLKS_ipd'event and RCLKS_ipd = '1') then

      case TO_X01(RBint_delayed) is
          when '1' =>
           null;
          when '0' =>

          if(RADDR < 0) then 
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          RPE_zd := 'X';
          if(TO_X01(RADDR0_delayed) = 'X') and (TO_X01(RADDR0_previous) /= 'X') then
             assert false
             report ": RADDR0 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR1_delayed) = 'X') and (TO_X01(RADDR1_previous) /= 'X') then
             assert false
             report ": RADDR1 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR2_delayed) = 'X') and (TO_X01(RADDR2_previous) /= 'X') then
             assert false
             report ": RADDR2 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR3_delayed) = 'X') and (TO_X01(RADDR3_previous) /= 'X') then
             assert false
             report ": RADDR3 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR4_delayed) = 'X') and (TO_X01(RADDR4_previous) /= 'X') then
             assert false
             report ": RADDR4 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR5_delayed) = 'X') and (TO_X01(RADDR5_previous) /= 'X') then
             assert false
             report ": RADDR5 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR6_delayed) = 'X') and (TO_X01(RADDR6_previous) /= 'X') then
             assert false
             report ": RADDR6 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR7_delayed) = 'X') and (TO_X01(RADDR7_previous) /= 'X') then
             assert false
             report ": RADDR7 unknown"
             severity Warning;
          end if;
          else  
            DO0_zd := memory_array(RADDR)(0);
            DO1_zd := memory_array(RADDR)(1);
            DO2_zd := memory_array(RADDR)(2);
            DO3_zd := memory_array(RADDR)(3);
            DO4_zd := memory_array(RADDR)(4);
            DO5_zd := memory_array(RADDR)(5);
            DO6_zd := memory_array(RADDR)(6);
            DO7_zd := memory_array(RADDR)(7);
            DO8_zd := memory_array(RADDR)(8);
            do_par  := DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR DO3_zd XOR DO2_zd XOR DO1_zd XOR DO0_zd;
            par_f <= do_par;
            if (do_par = 'X') then
              RPE_zd := 'X';
            elsif ( TO_X01 ( PARODD_delayed ) = 'X' ) then
              RPE_zd := 'X';
            else
              if (do_par /= PARODD_delayed) then
                RPE_zd  :=  '1';
              else
                RPE_zd  :=  '0';
              end if;
            end if;
        end if;

         when others =>
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          RPE_zd := 'X';
          if(TO_X01(RBint_previous) /= 'X') then
             assert false
             report ": RDB or RBLKB unknown "
             severity Warning;
           end if;
         end case;
       end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       RCLKS_previous  := RCLKS_ipd;
       RBint_previous := RBint_delayed;
       RBint_delayed  := RBint;
       WBint_previous  := WBint;
       RADDR0_previous := RADDR0_delayed;
       RADDR0_delayed  := RADDR0_ipd;
       RADDR1_previous := RADDR1_delayed;
       RADDR1_delayed  := RADDR1_ipd;
       RADDR2_previous := RADDR2_delayed;
       RADDR2_delayed  := RADDR2_ipd;
       RADDR3_previous := RADDR3_delayed;
       RADDR3_delayed  := RADDR3_ipd;
       RADDR4_previous := RADDR4_delayed;
       RADDR4_delayed  := RADDR4_ipd;
       RADDR5_previous := RADDR5_delayed;
       RADDR5_delayed  := RADDR5_ipd;
       RADDR6_previous := RADDR6_delayed;
       RADDR6_delayed  := RADDR6_ipd;
       RADDR7_previous := RADDR7_delayed;
       RADDR7_delayed  := RADDR7_ipd;
       WADDR0_previous := WADDR0_ipd;
       WADDR1_previous := WADDR1_ipd;
       WADDR2_previous := WADDR2_ipd;
       WADDR3_previous := WADDR3_ipd;
       WADDR4_previous := WADDR4_ipd;
       WADDR5_previous := WADDR5_ipd;
       WADDR6_previous := WADDR6_ipd;
       WADDR7_previous := WADDR7_ipd;
       PARODD_previous := PARODD_delayed; 
       PARODD_delayed  := PARODD_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
           OutSignal     => DOS,
           GlitchData    => DOS_GlitchData,
           OutSignalName => "DOS",
           OutTemp       => DOS_zd,
           Paths  =>  (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),
           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => WPE,
           GlitchData    => WPE_GlitchData,
           OutSignalName => "WPE",
           OutTemp       => WPE_zd,

           Paths  =>   (0 => (DI0_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI0_WPE),true),
                        1 => (DI1_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI1_WPE), true),
                        2 => (DI2_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI2_WPE), true),
                        3 => (DI3_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI3_WPE), true),
                        4 => (DI4_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI4_WPE), true),
                        5 => (DI5_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI5_WPE), true),
                        6 => (DI6_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI6_WPE), true),
                        7 => (DI7_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI7_WPE), true),
                        8 => (DI8_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI8_WPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => RPE,
           GlitchData    => RPE_GlitchData,
           OutSignalName => "RPE",
           OutTemp       => RPE_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_RPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
LIBRARY STD;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

USE std.textio.all;
USE ieee.std_logic_textio.all;
LIBRARY a500k;
USE a500k.all;

entity RAM256x9ASTP is 

   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                           : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                         : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                         : VitalDelayType := 0.000 ns;
 	tperiod_WRB                             : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WRB_RCLKS_negedge_posedge        : VitalDelayType := 0.000 ns;
 	thold_WRB_RCLKS_negedge_posedge         : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RCLKS_negedge_posedge      : VitalDelayType := 0.000 ns;
	thold_WBLKB_RCLKS_negedge_posedge       : VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');

ATTRIBUTE VITAL_LEVEL0 OF RAM256x9ASTP : entity IS True ;
END RAM256x9ASTP;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of RAM256x9ASTP is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal WADDR0_ipd : std_ulogic := 'X';
   signal WADDR1_ipd : std_ulogic := 'X';
   signal WADDR2_ipd : std_ulogic := 'X';
   signal WADDR3_ipd : std_ulogic := 'X';
   signal WADDR4_ipd : std_ulogic := 'X';
   signal WADDR5_ipd : std_ulogic := 'X';
   signal WADDR6_ipd : std_ulogic := 'X';
   signal WADDR7_ipd : std_ulogic := 'X';
   signal RADDR0_ipd : std_ulogic := 'X';
   signal RADDR1_ipd : std_ulogic := 'X';
   signal RADDR2_ipd : std_ulogic := 'X';
   signal RADDR3_ipd : std_ulogic := 'X';
   signal RADDR4_ipd : std_ulogic := 'X';
   signal RADDR5_ipd : std_ulogic := 'X';
   signal RADDR6_ipd : std_ulogic := 'X';
   signal RADDR7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

	-- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';
   signal INIT_MEM   : std_logic:= '0';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic:= 'X';
   signal par_f2     : std_logic:= 'X';

 begin  --  VITAL_ACT
   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (WADDR0_ipd, WADDR0, VitalExtendToFillDelay(tipd_WADDR0));
   VitalWireDelay (WADDR1_ipd, WADDR1, VitalExtendToFillDelay(tipd_WADDR1));
   VitalWireDelay (WADDR2_ipd, WADDR2, VitalExtendToFillDelay(tipd_WADDR2));
   VitalWireDelay (WADDR3_ipd, WADDR3, VitalExtendToFillDelay(tipd_WADDR3));
   VitalWireDelay (WADDR4_ipd, WADDR4, VitalExtendToFillDelay(tipd_WADDR4));
   VitalWireDelay (WADDR5_ipd, WADDR5, VitalExtendToFillDelay(tipd_WADDR5));
   VitalWireDelay (WADDR6_ipd, WADDR6, VitalExtendToFillDelay(tipd_WADDR6));
   VitalWireDelay (WADDR7_ipd, WADDR7, VitalExtendToFillDelay(tipd_WADDR7));
   VitalWireDelay (RADDR0_ipd, RADDR0, VitalExtendToFillDelay(tipd_RADDR0));
   VitalWireDelay (RADDR1_ipd, RADDR1, VitalExtendToFillDelay(tipd_RADDR1));
   VitalWireDelay (RADDR2_ipd, RADDR2, VitalExtendToFillDelay(tipd_RADDR2));
   VitalWireDelay (RADDR3_ipd, RADDR3, VitalExtendToFillDelay(tipd_RADDR3));
   VitalWireDelay (RADDR4_ipd, RADDR4, VitalExtendToFillDelay(tipd_RADDR4));
   VitalWireDelay (RADDR5_ipd, RADDR5, VitalExtendToFillDelay(tipd_RADDR5));
   VitalWireDelay (RADDR6_ipd, RADDR6, VitalExtendToFillDelay(tipd_RADDR6));
   VitalWireDelay (RADDR7_ipd, RADDR7, VitalExtendToFillDelay(tipd_RADDR7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

---------------------------------------------------------------
--                  Behavior Section                         --
---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);


    PROCESS
    BEGIN
      INIT_MEM <= '1';
      WAIT;
    END PROCESS;

    VITALBehavior : process (INIT_MEM, 
                          RADDR0_ipd, RADDR1_ipd, RADDR2_ipd, RADDR3_ipd, RADDR4_ipd, RADDR5_ipd, RADDR6_ipd, RADDR7_ipd, 
                          WADDR0_ipd, WADDR1_ipd, WADDR2_ipd, WADDR3_ipd, WADDR4_ipd, WADDR5_ipd, WADDR6_ipd, WADDR7_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd 
                          )

    -- some internal veriable declaration
     variable RAM_di_int         : std_logic_vector(8 downto 0);
     variable memory_array       : MEM_TYPE := (others =>(others => 'X'));
     variable do_par             : std_logic:= 'X';
     variable tmp_par            : std_logic:= 'X';
     variable tmp_par2           : std_logic:= 'X';
     variable wpe_var            : std_logic:= 'X';

     --  Read Timing Check Results
     variable Tviol_RADDR0_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR0_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR1_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR2_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR3_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR4_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR5_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR6_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR7_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable Tviol_WADDR0_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR0_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR0_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR0_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR0_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR1_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR1_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR1_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR1_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR2_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR2_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR2_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR2_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR3_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR3_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR3_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR3_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR4_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR4_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR4_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR4_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR5_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR5_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR5_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR5_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR6_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR6_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR6_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR6_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR7_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR7_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR7_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR7_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WRB_posedge      : X01                 := '0';
     variable TmDt_DI0_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI0_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WRB_posedge      : X01                 := '0';
     variable TmDt_DI1_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI1_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WRB_posedge      : X01                 := '0';
     variable TmDt_DI2_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI2_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WRB_posedge      : X01                 := '0';
     variable TmDt_DI3_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI3_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WRB_posedge      : X01                 := '0';
     variable TmDt_DI4_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI4_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WRB_posedge      : X01                 := '0';
     variable TmDt_DI5_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI5_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WRB_posedge      : X01                 := '0';
     variable TmDt_DI6_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI6_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WRB_posedge      : X01                 := '0';
     variable TmDt_DI7_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI7_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WRB_posedge      : X01                 := '0';
     variable TmDt_DI8_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI8_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WRB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WRB                  : X01                 := '0';
     variable PeriodData_WBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WBLKB                : X01                 := '0';
     variable Tviol_WRB_RCLKS_posedge    : X01 := '0';
     variable TmDt_WRB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_RCLKS_posedge  : X01 := '0';
     variable TmDt_WBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results

     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     variable DO0_zd : std_ulogic;
     variable DO1_zd : std_ulogic;
     variable DO2_zd : std_ulogic;
     variable DO3_zd : std_ulogic;
     variable DO4_zd : std_ulogic;
     variable DO5_zd : std_ulogic;
     variable DO6_zd : std_ulogic;
     variable DO7_zd : std_ulogic;
     variable DO8_zd : std_ulogic;
     variable RPE_zd : std_ulogic;
     variable WPE_zd : std_ulogic;
     variable DOS_zd : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData  : VitalGlitchDataType;
     variable DO1_GlitchData  : VitalGlitchDataType;
     variable DO2_GlitchData  : VitalGlitchDataType;
     variable DO3_GlitchData  : VitalGlitchDataType;
     variable DO4_GlitchData  : VitalGlitchDataType;
     variable DO5_GlitchData  : VitalGlitchDataType;
     variable DO6_GlitchData  : VitalGlitchDataType;
     variable DO7_GlitchData  : VitalGlitchDataType;
     variable DO8_GlitchData  : VitalGlitchDataType;
     variable DOS_GlitchData  : VitalGlitchDataType;

     -- last value variables
     variable RCLKS_previous  : std_ulogic := 'X';
     variable RBint_delayed   : std_ulogic := 'X';
     variable RBint_previous  : std_ulogic := 'X';
     variable WBint_previous  : std_ulogic := 'X';
     variable DIS_previous    : std_ulogic := 'X';
     variable RADDR0_delayed  : std_ulogic := 'X';
     variable RADDR1_delayed  : std_ulogic := 'X';
     variable RADDR2_delayed  : std_ulogic := 'X';
     variable RADDR3_delayed  : std_ulogic := 'X';
     variable RADDR4_delayed  : std_ulogic := 'X';
     variable RADDR5_delayed  : std_ulogic := 'X';
     variable RADDR6_delayed  : std_ulogic := 'X';
     variable RADDR7_delayed  : std_ulogic := 'X';
     variable RADDR0_previous : std_ulogic := 'X';
     variable RADDR1_previous : std_ulogic := 'X';
     variable RADDR2_previous : std_ulogic := 'X';
     variable RADDR3_previous : std_ulogic := 'X';
     variable RADDR4_previous : std_ulogic := 'X';
     variable RADDR5_previous : std_ulogic := 'X';
     variable RADDR6_previous : std_ulogic := 'X';
     variable RADDR7_previous : std_ulogic := 'X';
     variable WADDR0_previous : std_ulogic := 'X';
     variable WADDR1_previous : std_ulogic := 'X';
     variable WADDR2_previous : std_ulogic := 'X';
     variable WADDR3_previous : std_ulogic := 'X';
     variable WADDR4_previous : std_ulogic := 'X';
     variable WADDR5_previous : std_ulogic := 'X';
     variable WADDR6_previous : std_ulogic := 'X';
     variable WADDR7_previous : std_ulogic := 'X';

     variable PARODD_delayed  : std_ulogic := 'X';
     variable PARODD_previous : std_ulogic := 'X';
     variable Write_OK        : Boolean := FALSE;

     variable inline    : LINE;
     variable indata    : std_logic_vector(8 downto 0);
     variable resdata   : std_logic_vector(8 downto 0);
     variable i         : integer:=0;
     file     memfile   : text;
     variable status         : file_open_status;

 begin -- process VITALBehavior

  -----------------------------------------------------------
  --    Initialize memory file from MEMORYFILE string      --
  -----------------------------------------------------------

  if ( INIT_MEM'EVENT and INIT_MEM = '1') then
    file_open(status, memfile, MEMORYFILE, read_mode);
    if ( status=open_ok ) then
      while((i < 256) and (not ENDFILE(memfile))) loop
        readline(memfile,inline);
        read(inline,indata);
        resdata := indata;
        memory_array(i) := resdata;
        i := i+1;
      end loop;
    else
      assert ( MEMORYFILE'length = 0 )
        report "Failed to open RAM256x9ASTP memory initialization file in read mode"
        severity Note;
    end if;
    file_close(memfile);
  end if;


      WADDR := ((INT(WADDR7_ipd)*128)+(INT(WADDR6_ipd)*64)+(INT(
               WADDR5_ipd)*32) + (INT(WADDR4_ipd)*16) + 
               (INT(WADDR3_ipd)*8) + (INT(WADDR2_ipd)*4) + (INT(
               WADDR1_ipd)*2) + (INT(WADDR0_ipd)*1));
   -- Convert Read Address Signal to Integer
     if (RCLKS_ipd'EVENT AND RCLKS_ipd = '1') then
      RADDR := ((INT(RADDR7_delayed)*128)+(INT(RADDR6_delayed)*64)+(INT(
               RADDR5_delayed)*32) + (INT(RADDR4_delayed)*16) + 
               (INT(RADDR3_delayed)*8) + (INT(RADDR2_delayed)*4) + (INT(
               RADDR1_delayed)*2) + (INT(RADDR0_delayed)*1));
     end if;

if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

 -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9ASTP",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_negedge,
                             TmDt_WADDR0_WRB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR0_WRB_posedge_negedge,
                             tsetup_WADDR0_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_negedge,
                             TmDt_WADDR0_WRB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR0_WRB_negedge_negedge,
                             tsetup_WADDR0_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_negedge,
                             TmDt_WADDR1_WRB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR1_WRB_posedge_negedge,
                             tsetup_WADDR1_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_negedge,
                             TmDt_WADDR1_WRB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR1_WRB_negedge_negedge,
                             tsetup_WADDR1_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_negedge,
                             TmDt_WADDR2_WRB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR2_WRB_posedge_negedge,
                             tsetup_WADDR2_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_negedge,
                             TmDt_WADDR2_WRB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR2_WRB_negedge_negedge,
                             tsetup_WADDR2_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_negedge,
                             TmDt_WADDR3_WRB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR3_WRB_posedge_negedge,
                             tsetup_WADDR3_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_negedge,
                             TmDt_WADDR3_WRB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR3_WRB_negedge_negedge,
                             tsetup_WADDR3_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_negedge,
                             TmDt_WADDR4_WRB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR4_WRB_posedge_negedge,
                             tsetup_WADDR4_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_negedge,
                             TmDt_WADDR4_WRB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR4_WRB_negedge_negedge,
                             tsetup_WADDR4_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_negedge,
                             TmDt_WADDR5_WRB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR5_WRB_posedge_negedge,
                             tsetup_WADDR5_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_negedge,
                             TmDt_WADDR5_WRB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR5_WRB_negedge_negedge,
                             tsetup_WADDR5_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_negedge,
                             TmDt_WADDR6_WRB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR6_WRB_posedge_negedge,
                             tsetup_WADDR6_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_negedge,
                             TmDt_WADDR6_WRB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR6_WRB_negedge_negedge,
                             tsetup_WADDR6_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_negedge,
                             TmDt_WADDR7_WRB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR7_WRB_posedge_negedge,
                             tsetup_WADDR7_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_negedge,
                             TmDt_WADDR7_WRB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR7_WRB_negedge_negedge,
                             tsetup_WADDR7_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_negedge,
                             TmDt_WADDR0_WBLKB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR0_WBLKB_posedge_negedge,
                             tsetup_WADDR0_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_negedge,
                             TmDt_WADDR0_WBLKB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR0_WBLKB_negedge_negedge,
                             tsetup_WADDR0_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_negedge,
                             TmDt_WADDR1_WBLKB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR1_WBLKB_posedge_negedge,
                             tsetup_WADDR1_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_negedge,
                             TmDt_WADDR1_WBLKB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR1_WBLKB_negedge_negedge,
                             tsetup_WADDR1_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_negedge,
                             TmDt_WADDR2_WBLKB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR2_WBLKB_posedge_negedge,
                             tsetup_WADDR2_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_negedge,
                             TmDt_WADDR2_WBLKB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR2_WBLKB_negedge_negedge,
                             tsetup_WADDR2_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_negedge,
                             TmDt_WADDR3_WBLKB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR3_WBLKB_posedge_negedge,
                             tsetup_WADDR3_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_negedge,
                             TmDt_WADDR3_WBLKB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR3_WBLKB_negedge_negedge,
                             tsetup_WADDR3_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_negedge,
                             TmDt_WADDR4_WBLKB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR4_WBLKB_posedge_negedge,
                             tsetup_WADDR4_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_negedge,
                             TmDt_WADDR4_WBLKB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR4_WBLKB_negedge_negedge,
                             tsetup_WADDR4_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_negedge,
                             TmDt_WADDR5_WBLKB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR5_WBLKB_posedge_negedge,
                             tsetup_WADDR5_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_negedge,
                             TmDt_WADDR5_WBLKB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR5_WBLKB_negedge_negedge,
                             tsetup_WADDR5_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_negedge,
                             TmDt_WADDR6_WBLKB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR6_WBLKB_posedge_negedge,
                             tsetup_WADDR6_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_negedge,
                             TmDt_WADDR6_WBLKB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR6_WBLKB_negedge_negedge,
                             tsetup_WADDR6_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_negedge,
                             TmDt_WADDR7_WBLKB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR7_WBLKB_posedge_negedge,
                             tsetup_WADDR7_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_negedge,
                             TmDt_WADDR7_WBLKB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR7_WBLKB_negedge_negedge,
                             tsetup_WADDR7_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_posedge,
                             TmDt_WADDR0_WRB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WRB_posedge_posedge,
                             thold_WADDR0_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_posedge,
                             TmDt_WADDR0_WRB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WRB_negedge_posedge,
                             thold_WADDR0_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_posedge,
                             TmDt_WADDR1_WRB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WRB_posedge_posedge,
                             thold_WADDR1_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_posedge,
                             TmDt_WADDR1_WRB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WRB_negedge_posedge,
                             thold_WADDR1_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_posedge,
                             TmDt_WADDR2_WRB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WRB_posedge_posedge,
                             thold_WADDR2_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_posedge,
                             TmDt_WADDR2_WRB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WRB_negedge_posedge,
                             thold_WADDR2_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_posedge,
                             TmDt_WADDR3_WRB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WRB_posedge_posedge,
                             thold_WADDR3_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_posedge,
                             TmDt_WADDR3_WRB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WRB_negedge_posedge,
                             thold_WADDR3_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_posedge,
                             TmDt_WADDR4_WRB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WRB_posedge_posedge,
                             thold_WADDR4_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_posedge,
                             TmDt_WADDR4_WRB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WRB_negedge_posedge,
                             thold_WADDR4_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_posedge,
                             TmDt_WADDR5_WRB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WRB_posedge_posedge,
                             thold_WADDR5_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_posedge,
                             TmDt_WADDR5_WRB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WRB_negedge_posedge,
                             thold_WADDR5_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_posedge,
                             TmDt_WADDR6_WRB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WRB_posedge_posedge,
                             thold_WADDR6_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_posedge,
                             TmDt_WADDR6_WRB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WRB_negedge_posedge,
                             thold_WADDR6_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_posedge,
                             TmDt_WADDR7_WRB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WRB_posedge_posedge,
                             thold_WADDR7_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_posedge,
                             TmDt_WADDR7_WRB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WRB_negedge_posedge,
                             thold_WADDR7_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_posedge,
                             TmDt_WADDR0_WBLKB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WBLKB_posedge_posedge,
                             thold_WADDR0_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_posedge,
                             TmDt_WADDR0_WBLKB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WBLKB_negedge_posedge,
                             thold_WADDR0_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_posedge,
                             TmDt_WADDR1_WBLKB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WBLKB_posedge_posedge,
                             thold_WADDR1_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_posedge,
                             TmDt_WADDR1_WBLKB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WBLKB_negedge_posedge,
                             thold_WADDR1_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_posedge,
                             TmDt_WADDR2_WBLKB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WBLKB_posedge_posedge,
                             thold_WADDR2_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_posedge,
                             TmDt_WADDR2_WBLKB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WBLKB_negedge_posedge,
                             thold_WADDR2_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_posedge,
                             TmDt_WADDR3_WBLKB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WBLKB_posedge_posedge,
                             thold_WADDR3_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_posedge,
                             TmDt_WADDR3_WBLKB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WBLKB_negedge_posedge,
                             thold_WADDR3_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_posedge,
                             TmDt_WADDR4_WBLKB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WBLKB_posedge_posedge,
                             thold_WADDR4_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_posedge,
                             TmDt_WADDR4_WBLKB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WBLKB_negedge_posedge,
                             thold_WADDR4_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_posedge,
                             TmDt_WADDR5_WBLKB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WBLKB_posedge_posedge,
                             thold_WADDR5_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_posedge,
                             TmDt_WADDR5_WBLKB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WBLKB_negedge_posedge,
                             thold_WADDR5_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_posedge,
                             TmDt_WADDR6_WBLKB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WBLKB_posedge_posedge,
                             thold_WADDR6_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_posedge,
                             TmDt_WADDR6_WBLKB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WBLKB_negedge_posedge,
                             thold_WADDR6_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_posedge,
                             TmDt_WADDR7_WBLKB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WBLKB_posedge_posedge,
                             thold_WADDR7_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_posedge,
                             TmDt_WADDR7_WBLKB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WBLKB_negedge_posedge,
                             thold_WADDR7_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_posedge_posedge,
                             tsetup_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_negedge_posedge,
                             tsetup_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_posedge_posedge,
                             tsetup_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_negedge_posedge,
                             tsetup_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_posedge_posedge,
                             tsetup_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_negedge_posedge,
                             tsetup_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_posedge_posedge,
                             tsetup_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_negedge_posedge,
                             tsetup_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_posedge_posedge,
                             tsetup_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_negedge_posedge,
                             tsetup_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_posedge_posedge,
                             tsetup_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_negedge_posedge,
                             tsetup_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_posedge_posedge,
                             tsetup_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_negedge_posedge,
                             tsetup_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_posedge_posedge,
                             tsetup_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_negedge_posedge,
                             tsetup_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_posedge_posedge,
                             tsetup_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_negedge_posedge,
                             tsetup_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_posedge_posedge,
                             tsetup_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_negedge_posedge,
                             tsetup_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_posedge_posedge,
                             tsetup_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_negedge_posedge,
                             tsetup_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_posedge_posedge,
                             tsetup_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_negedge_posedge,
                             tsetup_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_posedge_posedge,
                             tsetup_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_negedge_posedge,
                             tsetup_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_posedge_posedge,
                             tsetup_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_negedge_posedge,
                             tsetup_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_posedge_posedge,
                             tsetup_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_negedge_posedge,
                             tsetup_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_posedge_posedge,
                             tsetup_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_negedge_posedge,
                             tsetup_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_posedge_posedge,
                             tsetup_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_negedge_posedge,
                             tsetup_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_posedge_posedge,
                             tsetup_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_negedge_posedge,
                             tsetup_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
      VitalPeriodPulseCheck ( Pviol_WBLKB,
                              PeriodData_WBLKB,
                              WBLKB_ipd, "WBLKB",
                              0.0 ns,
                              tperiod_WBLKB,
                              tpw_WBLKB_posedge,
                              tpw_WBLKB_negedge,
                              (To_X01(WRB_ipd) = '0'),
                              InstancePath & "/RAM256x9ASTP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_WRB,
                              PeriodData_WRB,
                              WRB_ipd, "WRB",
                              0.0 ns,
                              tperiod_WRB,
                              tpw_WRB_posedge,
                              tpw_WRB_negedge,
                              (To_X01(WBLKB_ipd) = '0'),
                              InstancePath & "/RAM256x9ASTP",
                              True,
                              True,
                              WARNING
                              );
   ------------------------------------------------------------
   --        Timing Checking for Read and write conflict     --
   ------------------------------------------------------------
       VitalSetupHoldCheck ( Tviol_WRB_RCLKS_posedge,
                             TmDt_WRB_RCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_WRB_RCLKS_negedge_posedge,
                             0.0 ns,
                             thold_WRB_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0') AND (To_X01(WBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_RCLKS_posedge,
                             TmDt_WBLKB_RCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_WBLKB_RCLKS_negedge_posedge,
                             0.0 ns,
                             thold_WBLKB_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0') AND (To_X01(WRB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

 end if;

   ------------------------------------------------------------
   --         WPE generating  block                            -
   ------------------------------------------------------------

      tmp_par  := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;
      if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
          ( TO_X01 ( DI7_ipd )    = 'X' ) or
          ( TO_X01 ( DI6_ipd )    = 'X' ) or
          ( TO_X01 ( DI5_ipd )    = 'X' ) or
          ( TO_X01 ( DI4_ipd )    = 'X' ) or
          ( TO_X01 ( DI3_ipd )    = 'X' ) or
          ( TO_X01 ( DI2_ipd )    = 'X' ) or
          ( TO_X01 ( DI1_ipd )    = 'X' ) or
          ( TO_X01 ( DI0_ipd )    = 'X' )
         ) then
        wpe_var  :=  'X';
      else
        if ( tmp_par /= PARODD_ipd ) then
          wpe_var  :=  '1';
        else
          wpe_var  :=  '0';
        end if;
      end if;
      RAM_di_int(8) := wpe_var;
      WPE_zd := wpe_var;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

    if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
    end if; 

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

   if (( TO_X01 ( WBint ) = '0' ) and ( TO_X01 ( WBint_previous ) = '1' )) then
     Write_OK := True;
   end if;


 -- async memory writing 
    if (TO_X01(WBint)='X') then
      if (TO_X01(WBint_previous) /= 'X') then
        assert false
        report ": WRB or WBLKB unknown"
        severity Warning;
      end if;
     elsif ( TO_X01(WBint) = '0' and Write_OK ) then
          if(WADDR < 0) then
           if((TO_X01(WADDR0_ipd) = 'X') and (TO_X01(WADDR0_previous) /= 'X')) then
             assert false
             report ": WADDR0 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR1_ipd) = 'X') and (TO_X01(WADDR1_previous) /= 'X')) then
             assert false
             report ": WADDR1 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR2_ipd) = 'X') and (TO_X01(WADDR2_previous) /= 'X')) then
             assert false
             report ": WADDR2 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR3_ipd) = 'X') and (TO_X01(WADDR3_previous) /= 'X')) then
             assert false
             report ": WADDR3 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR4_ipd) = 'X') and (TO_X01(WADDR4_previous) /= 'X')) then
             assert false
             report ": WADDR4 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR5_ipd) = 'X') and (TO_X01(WADDR5_previous) /= 'X')) then
             assert false
             report ": WADDR5 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR6_ipd) = 'X') and (TO_X01(WADDR6_previous) /= 'X')) then
             assert false
             report ": WADDR6 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR7_ipd) = 'X') and (TO_X01(WADDR7_previous) /= 'X')) then
             assert false
             report ": WADDR7 unknown, no data written ......"
             severity Warning;
           end if;
          else
             RAM_di_int(7 downto 0) :=DI7_ipd & DI6_ipd & DI5_ipd & DI4_ipd & DI3_ipd & DI2_ipd & DI1_ipd & DI0_ipd;
             memory_array(WADDR)  := RAM_di_int;
          end if;

    end if;


 -----------------------------------------------------------
 --  Read Functional Section                              --
 -----------------------------------------------------------


    if (TO_X01(RCLKS_ipd) = 'X') then
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          RPE_zd := 'X';
       if (TO_X01(RCLKS_previous) /= 'X') then
         assert false
         report ": RCLK unknown"
         severity Warning;
       end if;
    elsif(RCLKS_ipd'event and RCLKS_ipd = '1') then

      case TO_X01(RBint_delayed) is
          when '1' =>
           null;
          when '0' =>

          if(RADDR < 0) then 
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          if(TO_X01(RADDR0_delayed) = 'X') and (TO_X01(RADDR0_previous) /= 'X') then
             assert false
             report ": RADDR0 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR1_delayed) = 'X') and (TO_X01(RADDR1_previous) /= 'X') then
             assert false
             report ": RADDR1 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR2_delayed) = 'X') and (TO_X01(RADDR2_previous) /= 'X') then
             assert false
             report ": RADDR2 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR3_delayed) = 'X') and (TO_X01(RADDR3_previous) /= 'X') then
             assert false
             report ": RADDR3 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR4_delayed) = 'X') and (TO_X01(RADDR4_previous) /= 'X') then
             assert false
             report ": RADDR4 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR5_delayed) = 'X') and (TO_X01(RADDR5_previous) /= 'X') then
             assert false
             report ": RADDR5 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR6_delayed) = 'X') and (TO_X01(RADDR6_previous) /= 'X') then
             assert false
             report ": RADDR6 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR7_delayed) = 'X') and (TO_X01(RADDR7_previous) /= 'X') then
             assert false
             report ": RADDR7 unknown"
             severity Warning;
          end if;
          else  
            DO0_zd := memory_array(RADDR)(0);
            DO1_zd := memory_array(RADDR)(1);
            DO2_zd := memory_array(RADDR)(2);
            DO3_zd := memory_array(RADDR)(3);
            DO4_zd := memory_array(RADDR)(4);
            DO5_zd := memory_array(RADDR)(5);
            DO6_zd := memory_array(RADDR)(6);
            DO7_zd := memory_array(RADDR)(7);
            DO8_zd := memory_array(RADDR)(8);
        end if;

         when others =>
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          if(TO_X01(RBint_previous) /= 'X') then
             assert false
             report ": RDB or RBLKB unknown "
             severity Warning;
           end if;
         end case;
       end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       RCLKS_previous  := RCLKS_ipd;
       RBint_previous := RBint_delayed;
       RBint_delayed  := RBint;
       WBint_previous  := WBint;
       RADDR0_previous := RADDR0_delayed;
       RADDR0_delayed  := RADDR0_ipd;
       RADDR1_previous := RADDR1_delayed;
       RADDR1_delayed  := RADDR1_ipd;
       RADDR2_previous := RADDR2_delayed;
       RADDR2_delayed  := RADDR2_ipd;
       RADDR3_previous := RADDR3_delayed;
       RADDR3_delayed  := RADDR3_ipd;
       RADDR4_previous := RADDR4_delayed;
       RADDR4_delayed  := RADDR4_ipd;
       RADDR5_previous := RADDR5_delayed;
       RADDR5_delayed  := RADDR5_ipd;
       RADDR6_previous := RADDR6_delayed;
       RADDR6_delayed  := RADDR6_ipd;
       RADDR7_previous := RADDR7_delayed;
       RADDR7_delayed  := RADDR7_ipd;
       WADDR0_previous := WADDR0_ipd;
       WADDR1_previous := WADDR1_ipd;
       WADDR2_previous := WADDR2_ipd;
       WADDR3_previous := WADDR3_ipd;
       WADDR4_previous := WADDR4_ipd;
       WADDR5_previous := WADDR5_ipd;
       WADDR6_previous := WADDR6_ipd;
       WADDR7_previous := WADDR7_ipd;
       PARODD_previous := PARODD_delayed; 
       PARODD_delayed  := PARODD_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
           OutSignal     => DOS,
           GlitchData    => DOS_GlitchData,
           OutSignalName => "DOS",
           OutTemp       => DOS_zd,
           Paths  =>  (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),
           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
LIBRARY STD;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

USE std.textio.all;
USE ieee.std_logic_textio.all;
LIBRARY a500k;
USE a500k.all;

entity RAM256x9ASR is 

   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI0_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI1_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI2_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI3_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI4_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI5_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI6_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI7_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI8_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                           : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                         : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                         : VitalDelayType := 0.000 ns;
 	tperiod_WRB                             : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WRB_RCLKS_negedge_posedge        : VitalDelayType := 0.000 ns;
 	thold_WRB_RCLKS_negedge_posedge         : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RCLKS_negedge_posedge      : VitalDelayType := 0.000 ns;
	thold_WBLKB_RCLKS_negedge_posedge       : VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';
   WPE    :  OUT STD_LOGIC := 'X';
   RPE    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');

ATTRIBUTE VITAL_LEVEL0 OF RAM256x9ASR : entity IS True ;
END RAM256x9ASR;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of RAM256x9ASR is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal WADDR0_ipd : std_ulogic := 'X';
   signal WADDR1_ipd : std_ulogic := 'X';
   signal WADDR2_ipd : std_ulogic := 'X';
   signal WADDR3_ipd : std_ulogic := 'X';
   signal WADDR4_ipd : std_ulogic := 'X';
   signal WADDR5_ipd : std_ulogic := 'X';
   signal WADDR6_ipd : std_ulogic := 'X';
   signal WADDR7_ipd : std_ulogic := 'X';
   signal RADDR0_ipd : std_ulogic := 'X';
   signal RADDR1_ipd : std_ulogic := 'X';
   signal RADDR2_ipd : std_ulogic := 'X';
   signal RADDR3_ipd : std_ulogic := 'X';
   signal RADDR4_ipd : std_ulogic := 'X';
   signal RADDR5_ipd : std_ulogic := 'X';
   signal RADDR6_ipd : std_ulogic := 'X';
   signal RADDR7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

	-- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';
   signal INIT_MEM   : std_logic:= '0';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic:= 'X';
   signal par_f2     : std_logic:= 'X';

 begin  --  VITAL_ACT
   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (WADDR0_ipd, WADDR0, VitalExtendToFillDelay(tipd_WADDR0));
   VitalWireDelay (WADDR1_ipd, WADDR1, VitalExtendToFillDelay(tipd_WADDR1));
   VitalWireDelay (WADDR2_ipd, WADDR2, VitalExtendToFillDelay(tipd_WADDR2));
   VitalWireDelay (WADDR3_ipd, WADDR3, VitalExtendToFillDelay(tipd_WADDR3));
   VitalWireDelay (WADDR4_ipd, WADDR4, VitalExtendToFillDelay(tipd_WADDR4));
   VitalWireDelay (WADDR5_ipd, WADDR5, VitalExtendToFillDelay(tipd_WADDR5));
   VitalWireDelay (WADDR6_ipd, WADDR6, VitalExtendToFillDelay(tipd_WADDR6));
   VitalWireDelay (WADDR7_ipd, WADDR7, VitalExtendToFillDelay(tipd_WADDR7));
   VitalWireDelay (RADDR0_ipd, RADDR0, VitalExtendToFillDelay(tipd_RADDR0));
   VitalWireDelay (RADDR1_ipd, RADDR1, VitalExtendToFillDelay(tipd_RADDR1));
   VitalWireDelay (RADDR2_ipd, RADDR2, VitalExtendToFillDelay(tipd_RADDR2));
   VitalWireDelay (RADDR3_ipd, RADDR3, VitalExtendToFillDelay(tipd_RADDR3));
   VitalWireDelay (RADDR4_ipd, RADDR4, VitalExtendToFillDelay(tipd_RADDR4));
   VitalWireDelay (RADDR5_ipd, RADDR5, VitalExtendToFillDelay(tipd_RADDR5));
   VitalWireDelay (RADDR6_ipd, RADDR6, VitalExtendToFillDelay(tipd_RADDR6));
   VitalWireDelay (RADDR7_ipd, RADDR7, VitalExtendToFillDelay(tipd_RADDR7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

---------------------------------------------------------------
--                  Behavior Section                         --
---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);


    PROCESS
    BEGIN
      INIT_MEM <= '1';
      WAIT;
    END PROCESS;

    VITALBehavior : process (INIT_MEM, 
                          RADDR0_ipd, RADDR1_ipd, RADDR2_ipd, RADDR3_ipd, RADDR4_ipd, RADDR5_ipd, RADDR6_ipd, RADDR7_ipd, 
                          WADDR0_ipd, WADDR1_ipd, WADDR2_ipd, WADDR3_ipd, WADDR4_ipd, WADDR5_ipd, WADDR6_ipd, WADDR7_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd 
                          )

    -- some internal veriable declaration
     variable RAM_di_int         : std_logic_vector(8 downto 0);
     variable memory_array       : MEM_TYPE := (others =>(others => 'X'));
     variable do_par             : std_logic:= 'X';
     variable tmp_par            : std_logic:= 'X';
     variable tmp_par2           : std_logic:= 'X';
     variable wpe_var            : std_logic:= 'X';

     --  Read Timing Check Results
     variable Tviol_RADDR0_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR0_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR1_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR2_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR3_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR4_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR5_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR6_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR7_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable Tviol_WADDR0_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR0_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR0_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR0_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR0_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR1_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR1_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR1_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR1_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR2_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR2_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR2_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR2_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR3_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR3_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR3_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR3_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR4_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR4_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR4_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR4_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR5_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR5_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR5_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR5_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR6_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR6_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR6_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR6_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR7_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR7_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR7_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR7_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WRB_posedge      : X01                 := '0';
     variable TmDt_DI0_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI0_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WRB_posedge      : X01                 := '0';
     variable TmDt_DI1_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI1_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WRB_posedge      : X01                 := '0';
     variable TmDt_DI2_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI2_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WRB_posedge      : X01                 := '0';
     variable TmDt_DI3_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI3_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WRB_posedge      : X01                 := '0';
     variable TmDt_DI4_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI4_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WRB_posedge      : X01                 := '0';
     variable TmDt_DI5_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI5_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WRB_posedge      : X01                 := '0';
     variable TmDt_DI6_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI6_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WRB_posedge      : X01                 := '0';
     variable TmDt_DI7_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI7_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WRB_posedge      : X01                 := '0';
     variable TmDt_DI8_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI8_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WRB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WRB                  : X01                 := '0';
     variable PeriodData_WBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WBLKB                : X01                 := '0';
     variable Tviol_WRB_RCLKS_posedge    : X01 := '0';
     variable TmDt_WRB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_RCLKS_posedge  : X01 := '0';
     variable TmDt_WBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results

     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     variable DO0_zd : std_ulogic;
     variable DO1_zd : std_ulogic;
     variable DO2_zd : std_ulogic;
     variable DO3_zd : std_ulogic;
     variable DO4_zd : std_ulogic;
     variable DO5_zd : std_ulogic;
     variable DO6_zd : std_ulogic;
     variable DO7_zd : std_ulogic;
     variable DO8_zd : std_ulogic;
     variable RPE_zd : std_ulogic;
     variable WPE_zd : std_ulogic;
     variable DOS_zd : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData  : VitalGlitchDataType;
     variable DO1_GlitchData  : VitalGlitchDataType;
     variable DO2_GlitchData  : VitalGlitchDataType;
     variable DO3_GlitchData  : VitalGlitchDataType;
     variable DO4_GlitchData  : VitalGlitchDataType;
     variable DO5_GlitchData  : VitalGlitchDataType;
     variable DO6_GlitchData  : VitalGlitchDataType;
     variable DO7_GlitchData  : VitalGlitchDataType;
     variable DO8_GlitchData  : VitalGlitchDataType;
     variable RPE_GlitchData  : VitalGlitchDataType;
     variable WPE_GlitchData  : VitalGlitchDataType;
     variable DOS_GlitchData  : VitalGlitchDataType;

     -- last value variables
     variable RCLKS_previous  : std_ulogic := 'X';
     variable RBint_delayed   : std_ulogic := 'X';
     variable RBint_previous  : std_ulogic := 'X';
     variable WBint_previous  : std_ulogic := 'X';
     variable DIS_previous    : std_ulogic := 'X';
     variable RADDR0_delayed  : std_ulogic := 'X';
     variable RADDR1_delayed  : std_ulogic := 'X';
     variable RADDR2_delayed  : std_ulogic := 'X';
     variable RADDR3_delayed  : std_ulogic := 'X';
     variable RADDR4_delayed  : std_ulogic := 'X';
     variable RADDR5_delayed  : std_ulogic := 'X';
     variable RADDR6_delayed  : std_ulogic := 'X';
     variable RADDR7_delayed  : std_ulogic := 'X';
     variable RADDR0_previous : std_ulogic := 'X';
     variable RADDR1_previous : std_ulogic := 'X';
     variable RADDR2_previous : std_ulogic := 'X';
     variable RADDR3_previous : std_ulogic := 'X';
     variable RADDR4_previous : std_ulogic := 'X';
     variable RADDR5_previous : std_ulogic := 'X';
     variable RADDR6_previous : std_ulogic := 'X';
     variable RADDR7_previous : std_ulogic := 'X';
     variable WADDR0_previous : std_ulogic := 'X';
     variable WADDR1_previous : std_ulogic := 'X';
     variable WADDR2_previous : std_ulogic := 'X';
     variable WADDR3_previous : std_ulogic := 'X';
     variable WADDR4_previous : std_ulogic := 'X';
     variable WADDR5_previous : std_ulogic := 'X';
     variable WADDR6_previous : std_ulogic := 'X';
     variable WADDR7_previous : std_ulogic := 'X';

     --  Pipelined temporary results
     variable RPE_stg1        : std_ulogic := 'X';
     variable DO0_stg1        : std_ulogic := 'X';
     variable DO1_stg1        : std_ulogic := 'X';
     variable DO2_stg1        : std_ulogic := 'X';
     variable DO3_stg1        : std_ulogic := 'X';
     variable DO4_stg1        : std_ulogic := 'X';
     variable DO5_stg1        : std_ulogic := 'X';
     variable DO6_stg1        : std_ulogic := 'X';
     variable DO7_stg1        : std_ulogic := 'X';
     variable DO8_stg1        : std_ulogic := 'X';
 
     variable PARODD_delayed  : std_ulogic := 'X';
     variable PARODD_previous : std_ulogic := 'X';
     variable Write_OK        : Boolean := FALSE;
 
     variable inline    : LINE;
     variable indata    : std_logic_vector(8 downto 0);
     variable resdata   : std_logic_vector(8 downto 0);
     variable i         : integer:=0;
     file     memfile   : text;
     variable status         : file_open_status;

 begin -- process VITALBehavior

  -----------------------------------------------------------
  --    Initialize memory file from MEMORYFILE string      --
  -----------------------------------------------------------

  if ( INIT_MEM'EVENT and INIT_MEM = '1') then
    file_open(status, memfile, MEMORYFILE, read_mode);
    if ( status=open_ok ) then
      while((i < 256) and (not ENDFILE(memfile))) loop
        readline(memfile,inline);
        read(inline,indata);
        resdata := indata;
        memory_array(i) := resdata;
        i := i+1;
      end loop;
    else
      assert ( MEMORYFILE'length = 0 )
        report "Failed to open RAM256x9ASR memory initialization file in read mode"
        severity Note;
    end if;
    file_close(memfile);
  end if;


      WADDR := ((INT(WADDR7_ipd)*128)+(INT(WADDR6_ipd)*64)+(INT(
               WADDR5_ipd)*32) + (INT(WADDR4_ipd)*16) + 
               (INT(WADDR3_ipd)*8) + (INT(WADDR2_ipd)*4) + (INT(
               WADDR1_ipd)*2) + (INT(WADDR0_ipd)*1));
   -- Convert Read Address Signal to Integer
     if (RCLKS_ipd'EVENT AND RCLKS_ipd = '1') then
      RADDR := ((INT(RADDR7_delayed)*128)+(INT(RADDR6_delayed)*64)+(INT(
               RADDR5_delayed)*32) + (INT(RADDR4_delayed)*16) + 
               (INT(RADDR3_delayed)*8) + (INT(RADDR2_delayed)*4) + (INT(
               RADDR1_delayed)*2) + (INT(RADDR0_delayed)*1));
     end if;

if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

 -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9ASR",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_negedge,
                             TmDt_WADDR0_WRB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR0_WRB_posedge_negedge,
                             tsetup_WADDR0_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_negedge,
                             TmDt_WADDR0_WRB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR0_WRB_negedge_negedge,
                             tsetup_WADDR0_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_negedge,
                             TmDt_WADDR1_WRB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR1_WRB_posedge_negedge,
                             tsetup_WADDR1_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_negedge,
                             TmDt_WADDR1_WRB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR1_WRB_negedge_negedge,
                             tsetup_WADDR1_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_negedge,
                             TmDt_WADDR2_WRB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR2_WRB_posedge_negedge,
                             tsetup_WADDR2_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_negedge,
                             TmDt_WADDR2_WRB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR2_WRB_negedge_negedge,
                             tsetup_WADDR2_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_negedge,
                             TmDt_WADDR3_WRB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR3_WRB_posedge_negedge,
                             tsetup_WADDR3_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_negedge,
                             TmDt_WADDR3_WRB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR3_WRB_negedge_negedge,
                             tsetup_WADDR3_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_negedge,
                             TmDt_WADDR4_WRB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR4_WRB_posedge_negedge,
                             tsetup_WADDR4_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_negedge,
                             TmDt_WADDR4_WRB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR4_WRB_negedge_negedge,
                             tsetup_WADDR4_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_negedge,
                             TmDt_WADDR5_WRB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR5_WRB_posedge_negedge,
                             tsetup_WADDR5_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_negedge,
                             TmDt_WADDR5_WRB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR5_WRB_negedge_negedge,
                             tsetup_WADDR5_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_negedge,
                             TmDt_WADDR6_WRB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR6_WRB_posedge_negedge,
                             tsetup_WADDR6_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_negedge,
                             TmDt_WADDR6_WRB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR6_WRB_negedge_negedge,
                             tsetup_WADDR6_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_negedge,
                             TmDt_WADDR7_WRB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR7_WRB_posedge_negedge,
                             tsetup_WADDR7_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_negedge,
                             TmDt_WADDR7_WRB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR7_WRB_negedge_negedge,
                             tsetup_WADDR7_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_negedge,
                             TmDt_WADDR0_WBLKB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR0_WBLKB_posedge_negedge,
                             tsetup_WADDR0_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_negedge,
                             TmDt_WADDR0_WBLKB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR0_WBLKB_negedge_negedge,
                             tsetup_WADDR0_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_negedge,
                             TmDt_WADDR1_WBLKB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR1_WBLKB_posedge_negedge,
                             tsetup_WADDR1_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_negedge,
                             TmDt_WADDR1_WBLKB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR1_WBLKB_negedge_negedge,
                             tsetup_WADDR1_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_negedge,
                             TmDt_WADDR2_WBLKB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR2_WBLKB_posedge_negedge,
                             tsetup_WADDR2_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_negedge,
                             TmDt_WADDR2_WBLKB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR2_WBLKB_negedge_negedge,
                             tsetup_WADDR2_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_negedge,
                             TmDt_WADDR3_WBLKB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR3_WBLKB_posedge_negedge,
                             tsetup_WADDR3_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_negedge,
                             TmDt_WADDR3_WBLKB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR3_WBLKB_negedge_negedge,
                             tsetup_WADDR3_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_negedge,
                             TmDt_WADDR4_WBLKB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR4_WBLKB_posedge_negedge,
                             tsetup_WADDR4_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_negedge,
                             TmDt_WADDR4_WBLKB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR4_WBLKB_negedge_negedge,
                             tsetup_WADDR4_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_negedge,
                             TmDt_WADDR5_WBLKB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR5_WBLKB_posedge_negedge,
                             tsetup_WADDR5_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_negedge,
                             TmDt_WADDR5_WBLKB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR5_WBLKB_negedge_negedge,
                             tsetup_WADDR5_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_negedge,
                             TmDt_WADDR6_WBLKB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR6_WBLKB_posedge_negedge,
                             tsetup_WADDR6_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_negedge,
                             TmDt_WADDR6_WBLKB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR6_WBLKB_negedge_negedge,
                             tsetup_WADDR6_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_negedge,
                             TmDt_WADDR7_WBLKB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR7_WBLKB_posedge_negedge,
                             tsetup_WADDR7_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_negedge,
                             TmDt_WADDR7_WBLKB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR7_WBLKB_negedge_negedge,
                             tsetup_WADDR7_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_posedge,
                             TmDt_WADDR0_WRB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WRB_posedge_posedge,
                             thold_WADDR0_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_posedge,
                             TmDt_WADDR0_WRB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WRB_negedge_posedge,
                             thold_WADDR0_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_posedge,
                             TmDt_WADDR1_WRB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WRB_posedge_posedge,
                             thold_WADDR1_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_posedge,
                             TmDt_WADDR1_WRB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WRB_negedge_posedge,
                             thold_WADDR1_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_posedge,
                             TmDt_WADDR2_WRB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WRB_posedge_posedge,
                             thold_WADDR2_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_posedge,
                             TmDt_WADDR2_WRB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WRB_negedge_posedge,
                             thold_WADDR2_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_posedge,
                             TmDt_WADDR3_WRB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WRB_posedge_posedge,
                             thold_WADDR3_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_posedge,
                             TmDt_WADDR3_WRB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WRB_negedge_posedge,
                             thold_WADDR3_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_posedge,
                             TmDt_WADDR4_WRB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WRB_posedge_posedge,
                             thold_WADDR4_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_posedge,
                             TmDt_WADDR4_WRB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WRB_negedge_posedge,
                             thold_WADDR4_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_posedge,
                             TmDt_WADDR5_WRB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WRB_posedge_posedge,
                             thold_WADDR5_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_posedge,
                             TmDt_WADDR5_WRB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WRB_negedge_posedge,
                             thold_WADDR5_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_posedge,
                             TmDt_WADDR6_WRB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WRB_posedge_posedge,
                             thold_WADDR6_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_posedge,
                             TmDt_WADDR6_WRB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WRB_negedge_posedge,
                             thold_WADDR6_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_posedge,
                             TmDt_WADDR7_WRB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WRB_posedge_posedge,
                             thold_WADDR7_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_posedge,
                             TmDt_WADDR7_WRB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WRB_negedge_posedge,
                             thold_WADDR7_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_posedge,
                             TmDt_WADDR0_WBLKB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WBLKB_posedge_posedge,
                             thold_WADDR0_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_posedge,
                             TmDt_WADDR0_WBLKB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WBLKB_negedge_posedge,
                             thold_WADDR0_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_posedge,
                             TmDt_WADDR1_WBLKB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WBLKB_posedge_posedge,
                             thold_WADDR1_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_posedge,
                             TmDt_WADDR1_WBLKB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WBLKB_negedge_posedge,
                             thold_WADDR1_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_posedge,
                             TmDt_WADDR2_WBLKB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WBLKB_posedge_posedge,
                             thold_WADDR2_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_posedge,
                             TmDt_WADDR2_WBLKB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WBLKB_negedge_posedge,
                             thold_WADDR2_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_posedge,
                             TmDt_WADDR3_WBLKB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WBLKB_posedge_posedge,
                             thold_WADDR3_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_posedge,
                             TmDt_WADDR3_WBLKB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WBLKB_negedge_posedge,
                             thold_WADDR3_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_posedge,
                             TmDt_WADDR4_WBLKB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WBLKB_posedge_posedge,
                             thold_WADDR4_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_posedge,
                             TmDt_WADDR4_WBLKB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WBLKB_negedge_posedge,
                             thold_WADDR4_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_posedge,
                             TmDt_WADDR5_WBLKB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WBLKB_posedge_posedge,
                             thold_WADDR5_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_posedge,
                             TmDt_WADDR5_WBLKB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WBLKB_negedge_posedge,
                             thold_WADDR5_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_posedge,
                             TmDt_WADDR6_WBLKB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WBLKB_posedge_posedge,
                             thold_WADDR6_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_posedge,
                             TmDt_WADDR6_WBLKB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WBLKB_negedge_posedge,
                             thold_WADDR6_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_posedge,
                             TmDt_WADDR7_WBLKB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WBLKB_posedge_posedge,
                             thold_WADDR7_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_posedge,
                             TmDt_WADDR7_WBLKB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WBLKB_negedge_posedge,
                             thold_WADDR7_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_posedge_posedge,
                             tsetup_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_negedge_posedge,
                             tsetup_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_posedge_posedge,
                             tsetup_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_negedge_posedge,
                             tsetup_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_posedge_posedge,
                             tsetup_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_negedge_posedge,
                             tsetup_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_posedge_posedge,
                             tsetup_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_negedge_posedge,
                             tsetup_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_posedge_posedge,
                             tsetup_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_negedge_posedge,
                             tsetup_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_posedge_posedge,
                             tsetup_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_negedge_posedge,
                             tsetup_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_posedge_posedge,
                             tsetup_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_negedge_posedge,
                             tsetup_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_posedge_posedge,
                             tsetup_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_negedge_posedge,
                             tsetup_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_posedge_posedge,
                             tsetup_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_negedge_posedge,
                             tsetup_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_posedge_posedge,
                             tsetup_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_negedge_posedge,
                             tsetup_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_posedge_posedge,
                             tsetup_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_negedge_posedge,
                             tsetup_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_posedge_posedge,
                             tsetup_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_negedge_posedge,
                             tsetup_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_posedge_posedge,
                             tsetup_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_negedge_posedge,
                             tsetup_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_posedge_posedge,
                             tsetup_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_negedge_posedge,
                             tsetup_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_posedge_posedge,
                             tsetup_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_negedge_posedge,
                             tsetup_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_posedge_posedge,
                             tsetup_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_negedge_posedge,
                             tsetup_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_posedge_posedge,
                             tsetup_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_negedge_posedge,
                             tsetup_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_posedge_posedge,
                             tsetup_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_negedge_posedge,
                             tsetup_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );
      VitalPeriodPulseCheck ( Pviol_WBLKB,
                              PeriodData_WBLKB,
                              WBLKB_ipd, "WBLKB",
                              0.0 ns,
                              tperiod_WBLKB,
                              tpw_WBLKB_posedge,
                              tpw_WBLKB_negedge,
                              (To_X01(WRB_ipd) = '0'),
                              InstancePath & "/RAM256x9ASR",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_WRB,
                              PeriodData_WRB,
                              WRB_ipd, "WRB",
                              0.0 ns,
                              tperiod_WRB,
                              tpw_WRB_posedge,
                              tpw_WRB_negedge,
                              (To_X01(WBLKB_ipd) = '0'),
                              InstancePath & "/RAM256x9ASR",
                              True,
                              True,
                              WARNING
                              );
   ------------------------------------------------------------
   --        Timing Checking for Read and write conflict     --
   ------------------------------------------------------------
       VitalSetupHoldCheck ( Tviol_WRB_RCLKS_posedge,
                             TmDt_WRB_RCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_WRB_RCLKS_negedge_posedge,
                             0.0 ns,
                             thold_WRB_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0') AND (To_X01(WBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_RCLKS_posedge,
                             TmDt_WBLKB_RCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_WBLKB_RCLKS_negedge_posedge,
                             0.0 ns,
                             thold_WBLKB_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0') AND (To_X01(WRB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9ASR",
                             True,
                             True,
                             WARNING
                             );

 end if;

   ------------------------------------------------------------
   --    wpe output                                           -
   ------------------------------------------------------------

   if ( PARODD_ipd'EVENT ) then
     RPE_zd := not RPE_zd;
     RPE_stg1 := not RPE_stg1;
     WPE_zd := not WPE_zd;
   end if;

   ------------------------------------------------------------
   --         WPE checking  block                            -
   ------------------------------------------------------------

     tmp_par  := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;
     tmp_par2 := (tmp_par xor DI8_ipd);

      if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
          ( TO_X01 ( DI8_ipd )    = 'X' ) or
          ( TO_X01 ( DI7_ipd )    = 'X' ) or
          ( TO_X01 ( DI6_ipd )    = 'X' ) or
          ( TO_X01 ( DI5_ipd )    = 'X' ) or
          ( TO_X01 ( DI4_ipd )    = 'X' ) or
          ( TO_X01 ( DI3_ipd )    = 'X' ) or
          ( TO_X01 ( DI2_ipd )    = 'X' ) or
          ( TO_X01 ( DI1_ipd )    = 'X' ) or
          ( TO_X01 ( DI0_ipd )    = 'X' )
         ) then
        wpe_var  :=  'X';
      else
        if ( tmp_par2 /= PARODD_ipd ) then
          wpe_var  :=  '1';
        else
          wpe_var  :=  '0';
        end if;
      end if;
     RAM_di_int(8) := DI8_ipd;
     WPE_zd := wpe_var;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

    if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
    end if; 

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

   if (( TO_X01 ( WBint ) = '0' ) and ( TO_X01 ( WBint_previous ) = '1' )) then
     Write_OK := True;
   end if;


 -- async memory writing 
    if (TO_X01(WBint)='X') then
      if (TO_X01(WBint_previous) /= 'X') then
        assert false
        report ": WRB or WBLKB unknown"
        severity Warning;
      end if;
     elsif ( TO_X01(WBint) = '0' and Write_OK ) then
          if(WADDR < 0) then
           if((TO_X01(WADDR0_ipd) = 'X') and (TO_X01(WADDR0_previous) /= 'X')) then
             assert false
             report ": WADDR0 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR1_ipd) = 'X') and (TO_X01(WADDR1_previous) /= 'X')) then
             assert false
             report ": WADDR1 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR2_ipd) = 'X') and (TO_X01(WADDR2_previous) /= 'X')) then
             assert false
             report ": WADDR2 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR3_ipd) = 'X') and (TO_X01(WADDR3_previous) /= 'X')) then
             assert false
             report ": WADDR3 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR4_ipd) = 'X') and (TO_X01(WADDR4_previous) /= 'X')) then
             assert false
             report ": WADDR4 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR5_ipd) = 'X') and (TO_X01(WADDR5_previous) /= 'X')) then
             assert false
             report ": WADDR5 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR6_ipd) = 'X') and (TO_X01(WADDR6_previous) /= 'X')) then
             assert false
             report ": WADDR6 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR7_ipd) = 'X') and (TO_X01(WADDR7_previous) /= 'X')) then
             assert false
             report ": WADDR7 unknown, no data written ......"
             severity Warning;
           end if;
          else
             RAM_di_int(7 downto 0) :=DI7_ipd & DI6_ipd & DI5_ipd & DI4_ipd & DI3_ipd & DI2_ipd & DI1_ipd & DI0_ipd;
             memory_array(WADDR)  := RAM_di_int;
          end if;

    end if;


 -----------------------------------------------------------
 --  Read Functional Section                              --
 -----------------------------------------------------------


    if (TO_X01(RCLKS_ipd) = 'X') then
       DO0_stg1 := 'X';
       DO1_stg1 := 'X';
       DO2_stg1 := 'X';
       DO3_stg1 := 'X';
       DO4_stg1 := 'X';
       DO5_stg1 := 'X';
       DO6_stg1 := 'X';
       DO7_stg1 := 'X';
       DO8_stg1 := 'X';
       RPE_stg1 := 'X';
       if (TO_X01(RCLKS_previous) /= 'X') then
         assert false
         report ": RCLK unknown"
         severity Warning;
       end if;
    elsif(RCLKS_ipd'event and RCLKS_ipd = '1') then

      DO0_zd := DO0_stg1;
      DO1_zd := DO1_stg1;
      DO2_zd := DO2_stg1;
      DO3_zd := DO3_stg1;
      DO4_zd := DO4_stg1;
      DO5_zd := DO5_stg1;
      DO6_zd := DO6_stg1;
      DO7_zd := DO7_stg1;
      DO8_zd := DO8_stg1;
      RPE_zd := RPE_stg1;

      case TO_X01(RBint_delayed) is
          when '1' =>
           null;
          when '0' =>

          if(RADDR < 0) then 
          DO0_stg1 := 'X';
          DO1_stg1 := 'X';
          DO2_stg1 := 'X';
          DO3_stg1 := 'X';
          DO4_stg1 := 'X';
          DO5_stg1 := 'X';
          DO6_stg1 := 'X';
          DO7_stg1 := 'X';
          DO8_stg1 := 'X';
          RPE_stg1 := 'X';
          if(TO_X01(RADDR0_delayed) = 'X') and (TO_X01(RADDR0_previous) /= 'X') then
             assert false
             report ": RADDR0 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR1_delayed) = 'X') and (TO_X01(RADDR1_previous) /= 'X') then
             assert false
             report ": RADDR1 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR2_delayed) = 'X') and (TO_X01(RADDR2_previous) /= 'X') then
             assert false
             report ": RADDR2 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR3_delayed) = 'X') and (TO_X01(RADDR3_previous) /= 'X') then
             assert false
             report ": RADDR3 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR4_delayed) = 'X') and (TO_X01(RADDR4_previous) /= 'X') then
             assert false
             report ": RADDR4 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR5_delayed) = 'X') and (TO_X01(RADDR5_previous) /= 'X') then
             assert false
             report ": RADDR5 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR6_delayed) = 'X') and (TO_X01(RADDR6_previous) /= 'X') then
             assert false
             report ": RADDR6 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR7_delayed) = 'X') and (TO_X01(RADDR7_previous) /= 'X') then
             assert false
             report ": RADDR7 unknown"
             severity Warning;
          end if;
          else  
            DO0_stg1 :=memory_array(RADDR)(0);
            DO1_stg1 :=memory_array(RADDR)(1);
            DO2_stg1 :=memory_array(RADDR)(2);
            DO3_stg1 :=memory_array(RADDR)(3);
            DO4_stg1 :=memory_array(RADDR)(4);
            DO5_stg1 :=memory_array(RADDR)(5);
            DO6_stg1 :=memory_array(RADDR)(6);
            DO7_stg1 :=memory_array(RADDR)(7);
            DO8_stg1 :=memory_array(RADDR)(8);
            do_par  := DO8_stg1 XOR DO7_stg1 XOR DO6_stg1 XOR DO5_stg1 XOR DO4_stg1 XOR DO3_stg1 XOR DO2_stg1 XOR DO1_stg1 XOR DO0_stg1;
            par_f <= do_par;
            if ( do_par = 'X' ) then
              RPE_stg1 := 'X';
            elsif ( TO_X01 ( PARODD_delayed ) = 'X' ) then
              RPE_stg1 := 'X';
            else
              if ( do_par /= PARODD_delayed ) then
                RPE_stg1  :=  '1';
              else
                RPE_stg1  :=  '0';
              end if;
            end if;
        end if;

         when others =>
          DO0_stg1 := 'X';
          DO1_stg1 := 'X';
          DO2_stg1 := 'X';
          DO3_stg1 := 'X';
          DO4_stg1 := 'X';
          DO5_stg1 := 'X';
          DO6_stg1 := 'X';
          DO7_stg1 := 'X';
          DO8_stg1 := 'X';
          RPE_stg1 := 'X';
          if(TO_X01(RBint_previous) /= 'X') then
             assert false
             report ": RDB or RBLKB unknown "
             severity Warning;
           end if;
         end case;
       end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       RCLKS_previous  := RCLKS_ipd;
       RBint_previous := RBint_delayed;
       RBint_delayed  := RBint;
       WBint_previous  := WBint;
       RADDR0_previous := RADDR0_delayed;
       RADDR0_delayed  := RADDR0_ipd;
       RADDR1_previous := RADDR1_delayed;
       RADDR1_delayed  := RADDR1_ipd;
       RADDR2_previous := RADDR2_delayed;
       RADDR2_delayed  := RADDR2_ipd;
       RADDR3_previous := RADDR3_delayed;
       RADDR3_delayed  := RADDR3_ipd;
       RADDR4_previous := RADDR4_delayed;
       RADDR4_delayed  := RADDR4_ipd;
       RADDR5_previous := RADDR5_delayed;
       RADDR5_delayed  := RADDR5_ipd;
       RADDR6_previous := RADDR6_delayed;
       RADDR6_delayed  := RADDR6_ipd;
       RADDR7_previous := RADDR7_delayed;
       RADDR7_delayed  := RADDR7_ipd;
       WADDR0_previous := WADDR0_ipd;
       WADDR1_previous := WADDR1_ipd;
       WADDR2_previous := WADDR2_ipd;
       WADDR3_previous := WADDR3_ipd;
       WADDR4_previous := WADDR4_ipd;
       WADDR5_previous := WADDR5_ipd;
       WADDR6_previous := WADDR6_ipd;
       WADDR7_previous := WADDR7_ipd;
       PARODD_previous := PARODD_delayed; 
       PARODD_delayed  := PARODD_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
           OutSignal     => DOS,
           GlitchData    => DOS_GlitchData,
           OutSignalName => "DOS",
           OutTemp       => DOS_zd,
           Paths  =>  (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),
           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => WPE,
           GlitchData    => WPE_GlitchData,
           OutSignalName => "WPE",
           OutTemp       => WPE_zd,

           Paths  =>   (0 => (DI0_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI0_WPE),true),
                        1 => (DI1_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI1_WPE), true),
                        2 => (DI2_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI2_WPE), true),
                        3 => (DI3_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI3_WPE), true),
                        4 => (DI4_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI4_WPE), true),
                        5 => (DI5_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI5_WPE), true),
                        6 => (DI6_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI6_WPE), true),
                        7 => (DI7_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI7_WPE), true),
                        8 => (DI8_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI8_WPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => RPE,
           GlitchData    => RPE_GlitchData,
           OutSignalName => "RPE",
           OutTemp       => RPE_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_RPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
LIBRARY STD;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

USE std.textio.all;
USE ieee.std_logic_textio.all;
LIBRARY a500k;
USE a500k.all;

entity RAM256x9ASRP is 

   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_negedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_negedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WRB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WRB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                           : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                         : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                         : VitalDelayType := 0.000 ns;
 	tperiod_WRB                             : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WRB_RCLKS_negedge_posedge        : VitalDelayType := 0.000 ns;
 	thold_WRB_RCLKS_negedge_posedge         : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RCLKS_negedge_posedge      : VitalDelayType := 0.000 ns;
	thold_WBLKB_RCLKS_negedge_posedge       : VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');

ATTRIBUTE VITAL_LEVEL0 OF RAM256x9ASRP : entity IS True ;
END RAM256x9ASRP;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of RAM256x9ASRP is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal WADDR0_ipd : std_ulogic := 'X';
   signal WADDR1_ipd : std_ulogic := 'X';
   signal WADDR2_ipd : std_ulogic := 'X';
   signal WADDR3_ipd : std_ulogic := 'X';
   signal WADDR4_ipd : std_ulogic := 'X';
   signal WADDR5_ipd : std_ulogic := 'X';
   signal WADDR6_ipd : std_ulogic := 'X';
   signal WADDR7_ipd : std_ulogic := 'X';
   signal RADDR0_ipd : std_ulogic := 'X';
   signal RADDR1_ipd : std_ulogic := 'X';
   signal RADDR2_ipd : std_ulogic := 'X';
   signal RADDR3_ipd : std_ulogic := 'X';
   signal RADDR4_ipd : std_ulogic := 'X';
   signal RADDR5_ipd : std_ulogic := 'X';
   signal RADDR6_ipd : std_ulogic := 'X';
   signal RADDR7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

	-- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';
   signal INIT_MEM   : std_logic:= '0';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic:= 'X';
   signal par_f2     : std_logic:= 'X';

 begin  --  VITAL_ACT
   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (WADDR0_ipd, WADDR0, VitalExtendToFillDelay(tipd_WADDR0));
   VitalWireDelay (WADDR1_ipd, WADDR1, VitalExtendToFillDelay(tipd_WADDR1));
   VitalWireDelay (WADDR2_ipd, WADDR2, VitalExtendToFillDelay(tipd_WADDR2));
   VitalWireDelay (WADDR3_ipd, WADDR3, VitalExtendToFillDelay(tipd_WADDR3));
   VitalWireDelay (WADDR4_ipd, WADDR4, VitalExtendToFillDelay(tipd_WADDR4));
   VitalWireDelay (WADDR5_ipd, WADDR5, VitalExtendToFillDelay(tipd_WADDR5));
   VitalWireDelay (WADDR6_ipd, WADDR6, VitalExtendToFillDelay(tipd_WADDR6));
   VitalWireDelay (WADDR7_ipd, WADDR7, VitalExtendToFillDelay(tipd_WADDR7));
   VitalWireDelay (RADDR0_ipd, RADDR0, VitalExtendToFillDelay(tipd_RADDR0));
   VitalWireDelay (RADDR1_ipd, RADDR1, VitalExtendToFillDelay(tipd_RADDR1));
   VitalWireDelay (RADDR2_ipd, RADDR2, VitalExtendToFillDelay(tipd_RADDR2));
   VitalWireDelay (RADDR3_ipd, RADDR3, VitalExtendToFillDelay(tipd_RADDR3));
   VitalWireDelay (RADDR4_ipd, RADDR4, VitalExtendToFillDelay(tipd_RADDR4));
   VitalWireDelay (RADDR5_ipd, RADDR5, VitalExtendToFillDelay(tipd_RADDR5));
   VitalWireDelay (RADDR6_ipd, RADDR6, VitalExtendToFillDelay(tipd_RADDR6));
   VitalWireDelay (RADDR7_ipd, RADDR7, VitalExtendToFillDelay(tipd_RADDR7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

---------------------------------------------------------------
--                  Behavior Section                         --
---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);


    PROCESS
    BEGIN
      INIT_MEM <= '1';
      WAIT;
    END PROCESS;

    VITALBehavior : process (INIT_MEM, 
                          RADDR0_ipd, RADDR1_ipd, RADDR2_ipd, RADDR3_ipd, RADDR4_ipd, RADDR5_ipd, RADDR6_ipd, RADDR7_ipd, 
                          WADDR0_ipd, WADDR1_ipd, WADDR2_ipd, WADDR3_ipd, WADDR4_ipd, WADDR5_ipd, WADDR6_ipd, WADDR7_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd 
                          )

    -- some internal veriable declaration
     variable RAM_di_int         : std_logic_vector(8 downto 0);
     variable memory_array       : MEM_TYPE := (others =>(others => 'X'));
     variable do_par             : std_logic:= 'X';
     variable tmp_par            : std_logic:= 'X';
     variable tmp_par2           : std_logic:= 'X';
     variable wpe_var            : std_logic:= 'X';

     --  Read Timing Check Results
     variable Tviol_RADDR0_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR0_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR1_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR2_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR3_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR4_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR5_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR6_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR7_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable Tviol_WADDR0_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR0_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR0_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR0_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR0_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR0_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR1_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR1_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR1_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR1_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR2_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR2_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR2_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR2_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR3_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR3_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR3_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR3_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR4_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR4_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR4_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR4_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR5_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR5_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR5_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR5_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR6_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR6_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR6_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR6_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WRB_negedge   : X01                 := '0';
     variable TmDt_WADDR7_WRB_negedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WRB_posedge   : X01                 := '0';
     variable TmDt_WADDR7_WRB_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WBLKB_negedge : X01                 := '0';
     variable TmDt_WADDR7_WBLKB_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WBLKB_posedge : X01                 := '0';
     variable TmDt_WADDR7_WBLKB_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WRB_posedge      : X01                 := '0';
     variable TmDt_DI0_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI0_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WRB_posedge      : X01                 := '0';
     variable TmDt_DI1_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI1_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WRB_posedge      : X01                 := '0';
     variable TmDt_DI2_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI2_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WRB_posedge      : X01                 := '0';
     variable TmDt_DI3_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI3_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WRB_posedge      : X01                 := '0';
     variable TmDt_DI4_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI4_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WRB_posedge      : X01                 := '0';
     variable TmDt_DI5_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI5_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WRB_posedge      : X01                 := '0';
     variable TmDt_DI6_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI6_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WRB_posedge      : X01                 := '0';
     variable TmDt_DI7_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI7_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WRB_posedge      : X01                 := '0';
     variable TmDt_DI8_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI8_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WRB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WRB                  : X01                 := '0';
     variable PeriodData_WBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WBLKB                : X01                 := '0';
     variable Tviol_WRB_RCLKS_posedge    : X01 := '0';
     variable TmDt_WRB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_RCLKS_posedge  : X01 := '0';
     variable TmDt_WBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results

     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     variable DO0_zd : std_ulogic;
     variable DO1_zd : std_ulogic;
     variable DO2_zd : std_ulogic;
     variable DO3_zd : std_ulogic;
     variable DO4_zd : std_ulogic;
     variable DO5_zd : std_ulogic;
     variable DO6_zd : std_ulogic;
     variable DO7_zd : std_ulogic;
     variable DO8_zd : std_ulogic;
     variable RPE_zd : std_ulogic;
     variable WPE_zd : std_ulogic;
     variable DOS_zd : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData  : VitalGlitchDataType;
     variable DO1_GlitchData  : VitalGlitchDataType;
     variable DO2_GlitchData  : VitalGlitchDataType;
     variable DO3_GlitchData  : VitalGlitchDataType;
     variable DO4_GlitchData  : VitalGlitchDataType;
     variable DO5_GlitchData  : VitalGlitchDataType;
     variable DO6_GlitchData  : VitalGlitchDataType;
     variable DO7_GlitchData  : VitalGlitchDataType;
     variable DO8_GlitchData  : VitalGlitchDataType;
     variable DOS_GlitchData  : VitalGlitchDataType;

     -- last value variables
     variable RCLKS_previous  : std_ulogic := 'X';
     variable RBint_delayed   : std_ulogic := 'X';
     variable RBint_previous  : std_ulogic := 'X';
     variable WBint_previous  : std_ulogic := 'X';
     variable DIS_previous    : std_ulogic := 'X';
     variable RADDR0_delayed  : std_ulogic := 'X';
     variable RADDR1_delayed  : std_ulogic := 'X';
     variable RADDR2_delayed  : std_ulogic := 'X';
     variable RADDR3_delayed  : std_ulogic := 'X';
     variable RADDR4_delayed  : std_ulogic := 'X';
     variable RADDR5_delayed  : std_ulogic := 'X';
     variable RADDR6_delayed  : std_ulogic := 'X';
     variable RADDR7_delayed  : std_ulogic := 'X';
     variable RADDR0_previous : std_ulogic := 'X';
     variable RADDR1_previous : std_ulogic := 'X';
     variable RADDR2_previous : std_ulogic := 'X';
     variable RADDR3_previous : std_ulogic := 'X';
     variable RADDR4_previous : std_ulogic := 'X';
     variable RADDR5_previous : std_ulogic := 'X';
     variable RADDR6_previous : std_ulogic := 'X';
     variable RADDR7_previous : std_ulogic := 'X';
     variable WADDR0_previous : std_ulogic := 'X';
     variable WADDR1_previous : std_ulogic := 'X';
     variable WADDR2_previous : std_ulogic := 'X';
     variable WADDR3_previous : std_ulogic := 'X';
     variable WADDR4_previous : std_ulogic := 'X';
     variable WADDR5_previous : std_ulogic := 'X';
     variable WADDR6_previous : std_ulogic := 'X';
     variable WADDR7_previous : std_ulogic := 'X';

     --  Pipelined temporary results
     variable RPE_stg1        : std_ulogic := 'X';
     variable DO0_stg1        : std_ulogic := 'X';
     variable DO1_stg1        : std_ulogic := 'X';
     variable DO2_stg1        : std_ulogic := 'X';
     variable DO3_stg1        : std_ulogic := 'X';
     variable DO4_stg1        : std_ulogic := 'X';
     variable DO5_stg1        : std_ulogic := 'X';
     variable DO6_stg1        : std_ulogic := 'X';
     variable DO7_stg1        : std_ulogic := 'X';
     variable DO8_stg1        : std_ulogic := 'X';
 
     variable PARODD_delayed  : std_ulogic := 'X';
     variable PARODD_previous : std_ulogic := 'X';
     variable Write_OK        : Boolean := FALSE;
 
     variable inline    : LINE;
     variable indata    : std_logic_vector(8 downto 0);
     variable resdata   : std_logic_vector(8 downto 0);
     variable i         : integer:=0;
     file     memfile   : text;
     variable status         : file_open_status;
 
 begin -- process VITALBehavior

  -----------------------------------------------------------
  --    Initialize memory file from MEMORYFILE string      --
  -----------------------------------------------------------

  if ( INIT_MEM'EVENT and INIT_MEM = '1') then
    file_open(status, memfile, MEMORYFILE, read_mode);
    if ( status=open_ok ) then
      while((i < 256) and (not ENDFILE(memfile))) loop
        readline(memfile,inline);
        read(inline,indata);
        resdata := indata;
        memory_array(i) := resdata;
        i := i+1;
      end loop;
    else
      assert ( MEMORYFILE'length = 0 )
        report "Failed to open RAM256x9ASRP memory initialization file in read mode"
        severity Note;
    end if;
    file_close(memfile);
  end if;


      WADDR := ((INT(WADDR7_ipd)*128)+(INT(WADDR6_ipd)*64)+(INT(
               WADDR5_ipd)*32) + (INT(WADDR4_ipd)*16) + 
               (INT(WADDR3_ipd)*8) + (INT(WADDR2_ipd)*4) + (INT(
               WADDR1_ipd)*2) + (INT(WADDR0_ipd)*1));
   -- Convert Read Address Signal to Integer
     if (RCLKS_ipd'EVENT AND RCLKS_ipd = '1') then
      RADDR := ((INT(RADDR7_delayed)*128)+(INT(RADDR6_delayed)*64)+(INT(
               RADDR5_delayed)*32) + (INT(RADDR4_delayed)*16) + 
               (INT(RADDR3_delayed)*8) + (INT(RADDR2_delayed)*4) + (INT(
               RADDR1_delayed)*2) + (INT(RADDR0_delayed)*1));
     end if;

if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

 -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9ASRP",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_negedge,
                             TmDt_WADDR0_WRB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR0_WRB_posedge_negedge,
                             tsetup_WADDR0_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_negedge,
                             TmDt_WADDR0_WRB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR0_WRB_negedge_negedge,
                             tsetup_WADDR0_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_negedge,
                             TmDt_WADDR1_WRB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR1_WRB_posedge_negedge,
                             tsetup_WADDR1_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_negedge,
                             TmDt_WADDR1_WRB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR1_WRB_negedge_negedge,
                             tsetup_WADDR1_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_negedge,
                             TmDt_WADDR2_WRB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR2_WRB_posedge_negedge,
                             tsetup_WADDR2_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_negedge,
                             TmDt_WADDR2_WRB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR2_WRB_negedge_negedge,
                             tsetup_WADDR2_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_negedge,
                             TmDt_WADDR3_WRB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR3_WRB_posedge_negedge,
                             tsetup_WADDR3_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_negedge,
                             TmDt_WADDR3_WRB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR3_WRB_negedge_negedge,
                             tsetup_WADDR3_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_negedge,
                             TmDt_WADDR4_WRB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR4_WRB_posedge_negedge,
                             tsetup_WADDR4_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_negedge,
                             TmDt_WADDR4_WRB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR4_WRB_negedge_negedge,
                             tsetup_WADDR4_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_negedge,
                             TmDt_WADDR5_WRB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR5_WRB_posedge_negedge,
                             tsetup_WADDR5_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_negedge,
                             TmDt_WADDR5_WRB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR5_WRB_negedge_negedge,
                             tsetup_WADDR5_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_negedge,
                             TmDt_WADDR6_WRB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR6_WRB_posedge_negedge,
                             tsetup_WADDR6_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_negedge,
                             TmDt_WADDR6_WRB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR6_WRB_negedge_negedge,
                             tsetup_WADDR6_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_negedge,
                             TmDt_WADDR7_WRB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR7_WRB_posedge_negedge,
                             tsetup_WADDR7_WRB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_negedge,
                             TmDt_WADDR7_WRB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_WADDR7_WRB_negedge_negedge,
                             tsetup_WADDR7_WRB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBLKB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_negedge,
                             TmDt_WADDR0_WBLKB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR0_WBLKB_posedge_negedge,
                             tsetup_WADDR0_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_negedge,
                             TmDt_WADDR0_WBLKB_negedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR0_WBLKB_negedge_negedge,
                             tsetup_WADDR0_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_negedge,
                             TmDt_WADDR1_WBLKB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR1_WBLKB_posedge_negedge,
                             tsetup_WADDR1_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_negedge,
                             TmDt_WADDR1_WBLKB_negedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR1_WBLKB_negedge_negedge,
                             tsetup_WADDR1_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_negedge,
                             TmDt_WADDR2_WBLKB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR2_WBLKB_posedge_negedge,
                             tsetup_WADDR2_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_negedge,
                             TmDt_WADDR2_WBLKB_negedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR2_WBLKB_negedge_negedge,
                             tsetup_WADDR2_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_negedge,
                             TmDt_WADDR3_WBLKB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR3_WBLKB_posedge_negedge,
                             tsetup_WADDR3_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_negedge,
                             TmDt_WADDR3_WBLKB_negedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR3_WBLKB_negedge_negedge,
                             tsetup_WADDR3_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_negedge,
                             TmDt_WADDR4_WBLKB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR4_WBLKB_posedge_negedge,
                             tsetup_WADDR4_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_negedge,
                             TmDt_WADDR4_WBLKB_negedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR4_WBLKB_negedge_negedge,
                             tsetup_WADDR4_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_negedge,
                             TmDt_WADDR5_WBLKB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR5_WBLKB_posedge_negedge,
                             tsetup_WADDR5_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_negedge,
                             TmDt_WADDR5_WBLKB_negedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR5_WBLKB_negedge_negedge,
                             tsetup_WADDR5_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_negedge,
                             TmDt_WADDR6_WBLKB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR6_WBLKB_posedge_negedge,
                             tsetup_WADDR6_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_negedge,
                             TmDt_WADDR6_WBLKB_negedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR6_WBLKB_negedge_negedge,
                             tsetup_WADDR6_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_negedge,
                             TmDt_WADDR7_WBLKB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR7_WBLKB_posedge_negedge,
                             tsetup_WADDR7_WBLKB_posedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_negedge,
                             TmDt_WADDR7_WBLKB_negedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             tsetup_WADDR7_WBLKB_negedge_negedge,
                             tsetup_WADDR7_WBLKB_negedge_negedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WRB_ipd) = '0'),
                             '\',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_posedge,
                             TmDt_WADDR0_WRB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WRB_posedge_posedge,
                             thold_WADDR0_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WRB_posedge,
                             TmDt_WADDR0_WRB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WRB_negedge_posedge,
                             thold_WADDR0_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_posedge,
                             TmDt_WADDR1_WRB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WRB_posedge_posedge,
                             thold_WADDR1_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WRB_posedge,
                             TmDt_WADDR1_WRB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WRB_negedge_posedge,
                             thold_WADDR1_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_posedge,
                             TmDt_WADDR2_WRB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WRB_posedge_posedge,
                             thold_WADDR2_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WRB_posedge,
                             TmDt_WADDR2_WRB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WRB_negedge_posedge,
                             thold_WADDR2_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_posedge,
                             TmDt_WADDR3_WRB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WRB_posedge_posedge,
                             thold_WADDR3_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WRB_posedge,
                             TmDt_WADDR3_WRB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WRB_negedge_posedge,
                             thold_WADDR3_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_posedge,
                             TmDt_WADDR4_WRB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WRB_posedge_posedge,
                             thold_WADDR4_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WRB_posedge,
                             TmDt_WADDR4_WRB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WRB_negedge_posedge,
                             thold_WADDR4_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_posedge,
                             TmDt_WADDR5_WRB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WRB_posedge_posedge,
                             thold_WADDR5_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WRB_posedge,
                             TmDt_WADDR5_WRB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WRB_negedge_posedge,
                             thold_WADDR5_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_posedge,
                             TmDt_WADDR6_WRB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WRB_posedge_posedge,
                             thold_WADDR6_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WRB_posedge,
                             TmDt_WADDR6_WRB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WRB_negedge_posedge,
                             thold_WADDR6_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_posedge,
                             TmDt_WADDR7_WRB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WRB_posedge_posedge,
                             thold_WADDR7_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WRB_posedge,
                             TmDt_WADDR7_WRB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WRB_negedge_posedge,
                             thold_WADDR7_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_posedge,
                             TmDt_WADDR0_WBLKB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WBLKB_posedge_posedge,
                             thold_WADDR0_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR0_WBLKB_posedge,
                             TmDt_WADDR0_WBLKB_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR0_WBLKB_negedge_posedge,
                             thold_WADDR0_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_posedge,
                             TmDt_WADDR1_WBLKB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WBLKB_posedge_posedge,
                             thold_WADDR1_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR1_WBLKB_posedge,
                             TmDt_WADDR1_WBLKB_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR1_WBLKB_negedge_posedge,
                             thold_WADDR1_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_posedge,
                             TmDt_WADDR2_WBLKB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WBLKB_posedge_posedge,
                             thold_WADDR2_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR2_WBLKB_posedge,
                             TmDt_WADDR2_WBLKB_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR2_WBLKB_negedge_posedge,
                             thold_WADDR2_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_posedge,
                             TmDt_WADDR3_WBLKB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WBLKB_posedge_posedge,
                             thold_WADDR3_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR3_WBLKB_posedge,
                             TmDt_WADDR3_WBLKB_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR3_WBLKB_negedge_posedge,
                             thold_WADDR3_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_posedge,
                             TmDt_WADDR4_WBLKB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WBLKB_posedge_posedge,
                             thold_WADDR4_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR4_WBLKB_posedge,
                             TmDt_WADDR4_WBLKB_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR4_WBLKB_negedge_posedge,
                             thold_WADDR4_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_posedge,
                             TmDt_WADDR5_WBLKB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WBLKB_posedge_posedge,
                             thold_WADDR5_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR5_WBLKB_posedge,
                             TmDt_WADDR5_WBLKB_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR5_WBLKB_negedge_posedge,
                             thold_WADDR5_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_posedge,
                             TmDt_WADDR6_WBLKB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WBLKB_posedge_posedge,
                             thold_WADDR6_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR6_WBLKB_posedge,
                             TmDt_WADDR6_WBLKB_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR6_WBLKB_negedge_posedge,
                             thold_WADDR6_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_posedge,
                             TmDt_WADDR7_WBLKB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WBLKB_posedge_posedge,
                             thold_WADDR7_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_WADDR7_WBLKB_posedge,
                             TmDt_WADDR7_WBLKB_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_WADDR7_WBLKB_negedge_posedge,
                             thold_WADDR7_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_posedge_posedge,
                             tsetup_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_negedge_posedge,
                             tsetup_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_posedge_posedge,
                             tsetup_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_negedge_posedge,
                             tsetup_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_posedge_posedge,
                             tsetup_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_negedge_posedge,
                             tsetup_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_posedge_posedge,
                             tsetup_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_negedge_posedge,
                             tsetup_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_posedge_posedge,
                             tsetup_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_negedge_posedge,
                             tsetup_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_posedge_posedge,
                             tsetup_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_negedge_posedge,
                             tsetup_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_posedge_posedge,
                             tsetup_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_negedge_posedge,
                             tsetup_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_posedge_posedge,
                             tsetup_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_negedge_posedge,
                             tsetup_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_posedge_posedge,
                             tsetup_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_negedge_posedge,
                             tsetup_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_posedge_posedge,
                             tsetup_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_negedge_posedge,
                             tsetup_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_posedge_posedge,
                             tsetup_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_negedge_posedge,
                             tsetup_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_posedge_posedge,
                             tsetup_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_negedge_posedge,
                             tsetup_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_posedge_posedge,
                             tsetup_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_negedge_posedge,
                             tsetup_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_posedge_posedge,
                             tsetup_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_negedge_posedge,
                             tsetup_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_posedge_posedge,
                             tsetup_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_negedge_posedge,
                             tsetup_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_posedge_posedge,
                             tsetup_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_negedge_posedge,
                             tsetup_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_posedge_posedge,
                             tsetup_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_negedge_posedge,
                             tsetup_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_posedge_posedge,
                             tsetup_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_negedge_posedge,
                             tsetup_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
      VitalPeriodPulseCheck ( Pviol_WBLKB,
                              PeriodData_WBLKB,
                              WBLKB_ipd, "WBLKB",
                              0.0 ns,
                              tperiod_WBLKB,
                              tpw_WBLKB_posedge,
                              tpw_WBLKB_negedge,
                              (To_X01(WRB_ipd) = '0'),
                              InstancePath & "/RAM256x9ASRP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_WRB,
                              PeriodData_WRB,
                              WRB_ipd, "WRB",
                              0.0 ns,
                              tperiod_WRB,
                              tpw_WRB_posedge,
                              tpw_WRB_negedge,
                              (To_X01(WBLKB_ipd) = '0'),
                              InstancePath & "/RAM256x9ASRP",
                              True,
                              True,
                              WARNING
                              );
   ------------------------------------------------------------
   --        Timing Checking for Read and write conflict     --
   ------------------------------------------------------------
       VitalSetupHoldCheck ( Tviol_WRB_RCLKS_posedge,
                             TmDt_WRB_RCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_WRB_RCLKS_negedge_posedge,
                             0.0 ns,
                             thold_WRB_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0') AND (To_X01(WBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_RCLKS_posedge,
                             TmDt_WBLKB_RCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_WBLKB_RCLKS_negedge_posedge,
                             0.0 ns,
                             thold_WBLKB_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0') AND (To_X01(WRB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

 end if;

   ------------------------------------------------------------
   --         WPE generating  block                            -
   ------------------------------------------------------------

      tmp_par  := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;
      if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
          ( TO_X01 ( DI7_ipd )    = 'X' ) or
          ( TO_X01 ( DI6_ipd )    = 'X' ) or
          ( TO_X01 ( DI5_ipd )    = 'X' ) or
          ( TO_X01 ( DI4_ipd )    = 'X' ) or
          ( TO_X01 ( DI3_ipd )    = 'X' ) or
          ( TO_X01 ( DI2_ipd )    = 'X' ) or
          ( TO_X01 ( DI1_ipd )    = 'X' ) or
          ( TO_X01 ( DI0_ipd )    = 'X' )
         ) then
        wpe_var  :=  'X';
      else
        if ( tmp_par /= PARODD_ipd ) then
          wpe_var  :=  '1';
        else
          wpe_var  :=  '0';
        end if;
      end if;
      RAM_di_int(8) := wpe_var;
      WPE_zd := wpe_var;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

    if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
    end if; 

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

   if (( TO_X01 ( WBint ) = '0' ) and ( TO_X01 ( WBint_previous ) = '1' )) then
     Write_OK := True;
   end if;


 -- async memory writing 
    if (TO_X01(WBint)='X') then
      if (TO_X01(WBint_previous) /= 'X') then
        assert false
        report ": WRB or WBLKB unknown"
        severity Warning;
      end if;
     elsif ( TO_X01(WBint) = '0' and Write_OK ) then
          if(WADDR < 0) then
           if((TO_X01(WADDR0_ipd) = 'X') and (TO_X01(WADDR0_previous) /= 'X')) then
             assert false
             report ": WADDR0 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR1_ipd) = 'X') and (TO_X01(WADDR1_previous) /= 'X')) then
             assert false
             report ": WADDR1 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR2_ipd) = 'X') and (TO_X01(WADDR2_previous) /= 'X')) then
             assert false
             report ": WADDR2 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR3_ipd) = 'X') and (TO_X01(WADDR3_previous) /= 'X')) then
             assert false
             report ": WADDR3 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR4_ipd) = 'X') and (TO_X01(WADDR4_previous) /= 'X')) then
             assert false
             report ": WADDR4 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR5_ipd) = 'X') and (TO_X01(WADDR5_previous) /= 'X')) then
             assert false
             report ": WADDR5 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR6_ipd) = 'X') and (TO_X01(WADDR6_previous) /= 'X')) then
             assert false
             report ": WADDR6 unknown, no data written ......"
             severity Warning;
           end if;
           if((TO_X01(WADDR7_ipd) = 'X') and (TO_X01(WADDR7_previous) /= 'X')) then
             assert false
             report ": WADDR7 unknown, no data written ......"
             severity Warning;
           end if;
          else
             RAM_di_int(7 downto 0) :=DI7_ipd & DI6_ipd & DI5_ipd & DI4_ipd & DI3_ipd & DI2_ipd & DI1_ipd & DI0_ipd;
             memory_array(WADDR)  := RAM_di_int;
          end if;

    end if;


 -----------------------------------------------------------
 --  Read Functional Section                              --
 -----------------------------------------------------------


    if (TO_X01(RCLKS_ipd) = 'X') then
       DO0_stg1 := 'X';
       DO1_stg1 := 'X';
       DO2_stg1 := 'X';
       DO3_stg1 := 'X';
       DO4_stg1 := 'X';
       DO5_stg1 := 'X';
       DO6_stg1 := 'X';
       DO7_stg1 := 'X';
       DO8_stg1 := 'X';
       RPE_stg1 := 'X';
       if (TO_X01(RCLKS_previous) /= 'X') then
         assert false
         report ": RCLK unknown"
         severity Warning;
       end if;
    elsif(RCLKS_ipd'event and RCLKS_ipd = '1') then

      DO0_zd := DO0_stg1;
      DO1_zd := DO1_stg1;
      DO2_zd := DO2_stg1;
      DO3_zd := DO3_stg1;
      DO4_zd := DO4_stg1;
      DO5_zd := DO5_stg1;
      DO6_zd := DO6_stg1;
      DO7_zd := DO7_stg1;
      DO8_zd := DO8_stg1;
      RPE_zd := RPE_stg1;

      case TO_X01(RBint_delayed) is
          when '1' =>
           null;
          when '0' =>

          if(RADDR < 0) then 
          DO0_stg1 := 'X';
          DO1_stg1 := 'X';
          DO2_stg1 := 'X';
          DO3_stg1 := 'X';
          DO4_stg1 := 'X';
          DO5_stg1 := 'X';
          DO6_stg1 := 'X';
          DO7_stg1 := 'X';
          DO8_stg1 := 'X';
          if(TO_X01(RADDR0_delayed) = 'X') and (TO_X01(RADDR0_previous) /= 'X') then
             assert false
             report ": RADDR0 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR1_delayed) = 'X') and (TO_X01(RADDR1_previous) /= 'X') then
             assert false
             report ": RADDR1 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR2_delayed) = 'X') and (TO_X01(RADDR2_previous) /= 'X') then
             assert false
             report ": RADDR2 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR3_delayed) = 'X') and (TO_X01(RADDR3_previous) /= 'X') then
             assert false
             report ": RADDR3 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR4_delayed) = 'X') and (TO_X01(RADDR4_previous) /= 'X') then
             assert false
             report ": RADDR4 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR5_delayed) = 'X') and (TO_X01(RADDR5_previous) /= 'X') then
             assert false
             report ": RADDR5 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR6_delayed) = 'X') and (TO_X01(RADDR6_previous) /= 'X') then
             assert false
             report ": RADDR6 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR7_delayed) = 'X') and (TO_X01(RADDR7_previous) /= 'X') then
             assert false
             report ": RADDR7 unknown"
             severity Warning;
          end if;
          else  
            DO0_stg1 :=memory_array(RADDR)(0);
            DO1_stg1 :=memory_array(RADDR)(1);
            DO2_stg1 :=memory_array(RADDR)(2);
            DO3_stg1 :=memory_array(RADDR)(3);
            DO4_stg1 :=memory_array(RADDR)(4);
            DO5_stg1 :=memory_array(RADDR)(5);
            DO6_stg1 :=memory_array(RADDR)(6);
            DO7_stg1 :=memory_array(RADDR)(7);
            DO8_stg1 :=memory_array(RADDR)(8);
        end if;

         when others =>
          DO0_stg1 := 'X';
          DO1_stg1 := 'X';
          DO2_stg1 := 'X';
          DO3_stg1 := 'X';
          DO4_stg1 := 'X';
          DO5_stg1 := 'X';
          DO6_stg1 := 'X';
          DO7_stg1 := 'X';
          DO8_stg1 := 'X';
          if(TO_X01(RBint_previous) /= 'X') then
             assert false
             report ": RDB or RBLKB unknown "
             severity Warning;
           end if;
         end case;
       end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       RCLKS_previous  := RCLKS_ipd;
       RBint_previous := RBint_delayed;
       RBint_delayed  := RBint;
       WBint_previous  := WBint;
       RADDR0_previous := RADDR0_delayed;
       RADDR0_delayed  := RADDR0_ipd;
       RADDR1_previous := RADDR1_delayed;
       RADDR1_delayed  := RADDR1_ipd;
       RADDR2_previous := RADDR2_delayed;
       RADDR2_delayed  := RADDR2_ipd;
       RADDR3_previous := RADDR3_delayed;
       RADDR3_delayed  := RADDR3_ipd;
       RADDR4_previous := RADDR4_delayed;
       RADDR4_delayed  := RADDR4_ipd;
       RADDR5_previous := RADDR5_delayed;
       RADDR5_delayed  := RADDR5_ipd;
       RADDR6_previous := RADDR6_delayed;
       RADDR6_delayed  := RADDR6_ipd;
       RADDR7_previous := RADDR7_delayed;
       RADDR7_delayed  := RADDR7_ipd;
       WADDR0_previous := WADDR0_ipd;
       WADDR1_previous := WADDR1_ipd;
       WADDR2_previous := WADDR2_ipd;
       WADDR3_previous := WADDR3_ipd;
       WADDR4_previous := WADDR4_ipd;
       WADDR5_previous := WADDR5_ipd;
       WADDR6_previous := WADDR6_ipd;
       WADDR7_previous := WADDR7_ipd;
       PARODD_previous := PARODD_delayed; 
       PARODD_delayed  := PARODD_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
           OutSignal     => DOS,
           GlitchData    => DOS_GlitchData,
           OutSignalName => "DOS",
           OutTemp       => DOS_zd,
           Paths  =>  (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),
           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
LIBRARY STD;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

USE std.textio.all;
USE ieee.std_logic_textio.all;
LIBRARY a500k;
USE a500k.all;

entity RAM256x9SA is 

   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_WCLKS_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns,0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpw_RDB_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_RDB_negedge	        : VitalDelayType := 0.000 ns;
 	tperiod_RDB	        : VitalDelayType := 0.000 ns;
 	tpw_RBLKB_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RBLKB_negedge	: VitalDelayType := 0.000 ns;
 	tperiod_RBLKB	        : VitalDelayType := 0.000 ns;
 	tpw_RADDR0_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR0_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tpw_WCLKS_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                           : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_RDB_WCLKS_negedge_posedge       : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_WCLKS_negedge_posedge       : VitalDelayType := 0.000 ns;
 	tsetup_RADDR0_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR0_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR1_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR2_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR3_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR4_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR5_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR6_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR7_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	thold_RDB_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RBLKB_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR0_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR1_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR2_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR3_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR4_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR5_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR6_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR7_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';
   WPE    :  OUT STD_LOGIC := 'X';
   RPE    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   WCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');

ATTRIBUTE VITAL_LEVEL0 OF RAM256x9SA : entity IS True ;
END RAM256x9SA;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of RAM256x9SA is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal WADDR0_ipd : std_ulogic := 'X';
   signal WADDR1_ipd : std_ulogic := 'X';
   signal WADDR2_ipd : std_ulogic := 'X';
   signal WADDR3_ipd : std_ulogic := 'X';
   signal WADDR4_ipd : std_ulogic := 'X';
   signal WADDR5_ipd : std_ulogic := 'X';
   signal WADDR6_ipd : std_ulogic := 'X';
   signal WADDR7_ipd : std_ulogic := 'X';
   signal RADDR0_ipd : std_ulogic := 'X';
   signal RADDR1_ipd : std_ulogic := 'X';
   signal RADDR2_ipd : std_ulogic := 'X';
   signal RADDR3_ipd : std_ulogic := 'X';
   signal RADDR4_ipd : std_ulogic := 'X';
   signal RADDR5_ipd : std_ulogic := 'X';
   signal RADDR6_ipd : std_ulogic := 'X';
   signal RADDR7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal WCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

	-- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';
   signal INIT_MEM   : std_logic:= '0';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic:= 'X';
   signal par_f2     : std_logic:= 'X';

 begin  --  VITAL_ACT
   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (WADDR0_ipd, WADDR0, VitalExtendToFillDelay(tipd_WADDR0));
   VitalWireDelay (WADDR1_ipd, WADDR1, VitalExtendToFillDelay(tipd_WADDR1));
   VitalWireDelay (WADDR2_ipd, WADDR2, VitalExtendToFillDelay(tipd_WADDR2));
   VitalWireDelay (WADDR3_ipd, WADDR3, VitalExtendToFillDelay(tipd_WADDR3));
   VitalWireDelay (WADDR4_ipd, WADDR4, VitalExtendToFillDelay(tipd_WADDR4));
   VitalWireDelay (WADDR5_ipd, WADDR5, VitalExtendToFillDelay(tipd_WADDR5));
   VitalWireDelay (WADDR6_ipd, WADDR6, VitalExtendToFillDelay(tipd_WADDR6));
   VitalWireDelay (WADDR7_ipd, WADDR7, VitalExtendToFillDelay(tipd_WADDR7));
   VitalWireDelay (RADDR0_ipd, RADDR0, VitalExtendToFillDelay(tipd_RADDR0));
   VitalWireDelay (RADDR1_ipd, RADDR1, VitalExtendToFillDelay(tipd_RADDR1));
   VitalWireDelay (RADDR2_ipd, RADDR2, VitalExtendToFillDelay(tipd_RADDR2));
   VitalWireDelay (RADDR3_ipd, RADDR3, VitalExtendToFillDelay(tipd_RADDR3));
   VitalWireDelay (RADDR4_ipd, RADDR4, VitalExtendToFillDelay(tipd_RADDR4));
   VitalWireDelay (RADDR5_ipd, RADDR5, VitalExtendToFillDelay(tipd_RADDR5));
   VitalWireDelay (RADDR6_ipd, RADDR6, VitalExtendToFillDelay(tipd_RADDR6));
   VitalWireDelay (RADDR7_ipd, RADDR7, VitalExtendToFillDelay(tipd_RADDR7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (WCLKS_ipd, WCLKS, VitalExtendToFillDelay(tipd_WCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

---------------------------------------------------------------
--                  Behavior Section                         --
---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);


    PROCESS
    BEGIN
      INIT_MEM <= '1';
      WAIT;
    END PROCESS;

    VITALBehavior : process (INIT_MEM, 
                          RADDR0_ipd, RADDR1_ipd, RADDR2_ipd, RADDR3_ipd, RADDR4_ipd, RADDR5_ipd, RADDR6_ipd, RADDR7_ipd, 
                          WADDR0_ipd, WADDR1_ipd, WADDR2_ipd, WADDR3_ipd, WADDR4_ipd, WADDR5_ipd, WADDR6_ipd, WADDR7_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          WCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd 
                          )

    -- some internal veriable declaration
     variable RAM_di_int         : std_logic_vector(8 downto 0);
     variable memory_array       : MEM_TYPE := (others =>(others => 'X'));
     variable do_par             : std_logic:= 'X';
     variable tmp_par            : std_logic:= 'X';
     variable tmp_par2           : std_logic:= 'X';
     variable wpe_var            : std_logic:= 'X';

     --  Read Timing Check Results
     variable PeriodData_RDB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RDB                  : X01                 := '0';
     variable PeriodData_RBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RBLKB                : X01                  := '0';
     variable PeriodData_RADDR0          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR0               : X01                 := '0';
     variable PeriodData_RADDR1          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR1               : X01                 := '0';
     variable PeriodData_RADDR2          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR2               : X01                 := '0';
     variable PeriodData_RADDR3          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR3               : X01                 := '0';
     variable PeriodData_RADDR4          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR4               : X01                 := '0';
     variable PeriodData_RADDR5          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR5               : X01                 := '0';
     variable PeriodData_RADDR6          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR6               : X01                 := '0';
     variable PeriodData_RADDR7          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR7               : X01                 := '0';
     variable Tviol_WADDR0_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR0_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR1_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR2_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR3_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR4_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR5_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR6_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR7_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI0_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI1_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI2_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI3_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI4_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI5_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI6_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI7_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI8_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_WCLKS_posedge    : X01                 := '0';
     variable TmDt_WRB_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_WCLKS_posedge  : X01                 := '0';
     variable TmDt_WBLKB_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WCLKS                : X01                 := '0';
     variable Tviol_RDB_WCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_WCLKS_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_WCLKS_negedge    : X01                 := '0';
     variable TmDt_RDB_WCLKS_negedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_WCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_WCLKS_negedge  : X01                 := '0';
     variable TmDt_RBLKB_WCLKS_negedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR0_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR0_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR0_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR0_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR1_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR1_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR2_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR2_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR3_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR3_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR4_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR4_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR5_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR5_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR6_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR6_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR7_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR7_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results

     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     variable DO0_zd : std_ulogic;
     variable DO1_zd : std_ulogic;
     variable DO2_zd : std_ulogic;
     variable DO3_zd : std_ulogic;
     variable DO4_zd : std_ulogic;
     variable DO5_zd : std_ulogic;
     variable DO6_zd : std_ulogic;
     variable DO7_zd : std_ulogic;
     variable DO8_zd : std_ulogic;
     variable RPE_zd : std_ulogic;
     variable WPE_zd : std_ulogic;
     variable DOS_zd : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData  : VitalGlitchDataType;
     variable DO1_GlitchData  : VitalGlitchDataType;
     variable DO2_GlitchData  : VitalGlitchDataType;
     variable DO3_GlitchData  : VitalGlitchDataType;
     variable DO4_GlitchData  : VitalGlitchDataType;
     variable DO5_GlitchData  : VitalGlitchDataType;
     variable DO6_GlitchData  : VitalGlitchDataType;
     variable DO7_GlitchData  : VitalGlitchDataType;
     variable DO8_GlitchData  : VitalGlitchDataType;
     variable RPE_GlitchData  : VitalGlitchDataType;
     variable WPE_GlitchData  : VitalGlitchDataType;
     variable DOS_GlitchData  : VitalGlitchDataType;

     -- last value variables
     variable WCLKS_previous  : std_ulogic := 'X';
     variable RBint_previous  : std_ulogic := 'X';
     variable WBint_delayed   : std_ulogic := 'X';
     variable WBint_previous  : std_ulogic := 'X';
     variable DIS_previous    : std_ulogic := 'X';
     variable DI0_delayed     : std_ulogic := 'X';
     variable DI1_delayed     : std_ulogic := 'X';
     variable DI2_delayed     : std_ulogic := 'X';
     variable DI3_delayed     : std_ulogic := 'X';
     variable DI4_delayed     : std_ulogic := 'X';
     variable DI5_delayed     : std_ulogic := 'X';
     variable DI6_delayed     : std_ulogic := 'X';
     variable DI7_delayed     : std_ulogic := 'X';
     variable DI8_delayed     : std_ulogic := 'X';
     variable RADDR0_previous : std_ulogic := 'X';
     variable RADDR1_previous : std_ulogic := 'X';
     variable RADDR2_previous : std_ulogic := 'X';
     variable RADDR3_previous : std_ulogic := 'X';
     variable RADDR4_previous : std_ulogic := 'X';
     variable RADDR5_previous : std_ulogic := 'X';
     variable RADDR6_previous : std_ulogic := 'X';
     variable RADDR7_previous : std_ulogic := 'X';
     variable WADDR0_delayed  : std_ulogic := 'X';
     variable WADDR1_delayed  : std_ulogic := 'X';
     variable WADDR2_delayed  : std_ulogic := 'X';
     variable WADDR3_delayed  : std_ulogic := 'X';
     variable WADDR4_delayed  : std_ulogic := 'X';
     variable WADDR5_delayed  : std_ulogic := 'X';
     variable WADDR6_delayed  : std_ulogic := 'X';
     variable WADDR7_delayed  : std_ulogic := 'X';
     variable WADDR0_previous : std_ulogic := 'X';
     variable WADDR1_previous : std_ulogic := 'X';
     variable WADDR2_previous : std_ulogic := 'X';
     variable WADDR3_previous : std_ulogic := 'X';
     variable WADDR4_previous : std_ulogic := 'X';
     variable WADDR5_previous : std_ulogic := 'X';
     variable WADDR6_previous : std_ulogic := 'X';
     variable WADDR7_previous : std_ulogic := 'X';

     variable PARODD_delayed  : std_ulogic := 'X';
     variable PARODD_previous : std_ulogic := 'X';
 
     variable inline    : LINE;
     variable indata    : std_logic_vector(8 downto 0);
     variable resdata   : std_logic_vector(8 downto 0);
     variable i         : integer:=0;
     file     memfile   : text;
     variable status         : file_open_status;

 begin -- process VITALBehavior

  -----------------------------------------------------------
  --    Initialize memory file from MEMORYFILE string      --
  -----------------------------------------------------------


  if ( INIT_MEM'EVENT and INIT_MEM = '1') then
    file_open(status, memfile, MEMORYFILE, read_mode);
    if ( status=open_ok ) then
      while((i < 256) and (not ENDFILE(memfile))) loop
        readline(memfile,inline);
        read(inline,indata);
        resdata := indata;
        memory_array(i) := resdata;
        i := i+1;
      end loop;
    else
      assert ( MEMORYFILE'length = 0 )
        report "Failed to open RAM256x9SA memory initialization file in read mode"
        severity Note;
    end if;
    file_close(memfile);
  end if;


     if (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      WADDR := ((INT(WADDR7_delayed)*128)+(INT(WADDR6_delayed)*64)+(INT(
               WADDR5_delayed)*32) + (INT(WADDR4_delayed)*16) + 
               (INT(WADDR3_delayed)*8) + (INT(WADDR2_delayed)*4) + (INT(
               WADDR1_delayed)*2) + (INT(WADDR0_delayed)*1));
     end if;

   -- Convert Read Address Signal to Integer

      RADDR := ((INT(RADDR7_ipd)*128)+(INT(RADDR6_ipd)*64)+(INT(
               RADDR5_ipd)*32) + (INT(RADDR4_ipd)*16) + 
               (INT(RADDR3_ipd)*8) + (INT(RADDR2_ipd)*4) + (INT(
               RADDR1_ipd)*2) + (INT(RADDR0_ipd)*1));

if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

      VitalPeriodPulseCheck ( Pviol_RDB,
                              PeriodData_RDB,
                              RDB_ipd, "RDB",
                              0.0 ns,
                              tperiod_RDB,
                              tpw_RDB_posedge,
                              tpw_RDB_negedge,
                              (To_X01(RBLKB_ipd) = '0'),
                             InstancePath &"/RAM256x9SA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RBLKB,
                              PeriodData_RBLKB,
                              RBLKB_ipd, "RBLKB",
                              0.0 ns,
                              tperiod_RBLKB,
                              tpw_RBLKB_posedge,
                              tpw_RBLKB_negedge,
                              (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR0,
                              PeriodData_RADDR0,
                              RADDR0_ipd, "RADDR0",
                              0.0 ns,
                              tpw_RADDR0_posedge + tpw_RADDR0_posedge,
                              tpw_RADDR0_posedge,
                              tpw_RADDR0_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR1,
                              PeriodData_RADDR1,
                              RADDR1_ipd, "RADDR1",
                              0.0 ns,
                              tpw_RADDR1_posedge + tpw_RADDR1_posedge,
                              tpw_RADDR1_posedge,
                              tpw_RADDR1_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR2,
                              PeriodData_RADDR2,
                              RADDR2_ipd, "RADDR2",
                              0.0 ns,
                              tpw_RADDR2_posedge + tpw_RADDR2_posedge,
                              tpw_RADDR2_posedge,
                              tpw_RADDR2_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR3,
                              PeriodData_RADDR3,
                              RADDR3_ipd, "RADDR3",
                              0.0 ns,
                              tpw_RADDR3_posedge + tpw_RADDR3_posedge,
                              tpw_RADDR3_posedge,
                              tpw_RADDR3_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR4,
                              PeriodData_RADDR4,
                              RADDR4_ipd, "RADDR4",
                              0.0 ns,
                              tpw_RADDR4_posedge + tpw_RADDR4_posedge,
                              tpw_RADDR4_posedge,
                              tpw_RADDR4_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR5,
                              PeriodData_RADDR5,
                              RADDR5_ipd, "RADDR5",
                              0.0 ns,
                              tpw_RADDR5_posedge + tpw_RADDR5_posedge,
                              tpw_RADDR5_posedge,
                              tpw_RADDR5_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR6,
                              PeriodData_RADDR6,
                              RADDR6_ipd, "RADDR6",
                              0.0 ns,
                              tpw_RADDR6_posedge + tpw_RADDR6_posedge,
                              tpw_RADDR6_posedge,
                              tpw_RADDR6_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR7,
                              PeriodData_RADDR7,
                              RADDR7_ipd, "RADDR7",
                              0.0 ns,
                              tpw_RADDR7_posedge + tpw_RADDR7_posedge,
                              tpw_RADDR7_posedge,
                              tpw_RADDR7_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SA",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_WADDR0_WCLKS_posedge,
                             TmDt_WADDR0_WCLKS_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR0_WCLKS_posedge_posedge,
                             tsetup_WADDR0_WCLKS_posedge_posedge,
                             thold_WADDR0_WCLKS_posedge_posedge,
                             thold_WADDR0_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WCLKS_posedge,
                             TmDt_WADDR0_WCLKS_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR0_WCLKS_negedge_posedge,
                             tsetup_WADDR0_WCLKS_negedge_posedge,
                             thold_WADDR0_WCLKS_negedge_posedge,
                             thold_WADDR0_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WCLKS_posedge,
                             TmDt_WADDR1_WCLKS_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR1_WCLKS_posedge_posedge,
                             tsetup_WADDR1_WCLKS_posedge_posedge,
                             thold_WADDR1_WCLKS_posedge_posedge,
                             thold_WADDR1_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WCLKS_posedge,
                             TmDt_WADDR1_WCLKS_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR1_WCLKS_negedge_posedge,
                             tsetup_WADDR1_WCLKS_negedge_posedge,
                             thold_WADDR1_WCLKS_negedge_posedge,
                             thold_WADDR1_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WCLKS_posedge,
                             TmDt_WADDR2_WCLKS_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR2_WCLKS_posedge_posedge,
                             tsetup_WADDR2_WCLKS_posedge_posedge,
                             thold_WADDR2_WCLKS_posedge_posedge,
                             thold_WADDR2_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WCLKS_posedge,
                             TmDt_WADDR2_WCLKS_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR2_WCLKS_negedge_posedge,
                             tsetup_WADDR2_WCLKS_negedge_posedge,
                             thold_WADDR2_WCLKS_negedge_posedge,
                             thold_WADDR2_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WCLKS_posedge,
                             TmDt_WADDR3_WCLKS_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR3_WCLKS_posedge_posedge,
                             tsetup_WADDR3_WCLKS_posedge_posedge,
                             thold_WADDR3_WCLKS_posedge_posedge,
                             thold_WADDR3_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WCLKS_posedge,
                             TmDt_WADDR3_WCLKS_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR3_WCLKS_negedge_posedge,
                             tsetup_WADDR3_WCLKS_negedge_posedge,
                             thold_WADDR3_WCLKS_negedge_posedge,
                             thold_WADDR3_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WCLKS_posedge,
                             TmDt_WADDR4_WCLKS_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR4_WCLKS_posedge_posedge,
                             tsetup_WADDR4_WCLKS_posedge_posedge,
                             thold_WADDR4_WCLKS_posedge_posedge,
                             thold_WADDR4_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WCLKS_posedge,
                             TmDt_WADDR4_WCLKS_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR4_WCLKS_negedge_posedge,
                             tsetup_WADDR4_WCLKS_negedge_posedge,
                             thold_WADDR4_WCLKS_negedge_posedge,
                             thold_WADDR4_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WCLKS_posedge,
                             TmDt_WADDR5_WCLKS_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR5_WCLKS_posedge_posedge,
                             tsetup_WADDR5_WCLKS_posedge_posedge,
                             thold_WADDR5_WCLKS_posedge_posedge,
                             thold_WADDR5_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WCLKS_posedge,
                             TmDt_WADDR5_WCLKS_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR5_WCLKS_negedge_posedge,
                             tsetup_WADDR5_WCLKS_negedge_posedge,
                             thold_WADDR5_WCLKS_negedge_posedge,
                             thold_WADDR5_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WCLKS_posedge,
                             TmDt_WADDR6_WCLKS_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR6_WCLKS_posedge_posedge,
                             tsetup_WADDR6_WCLKS_posedge_posedge,
                             thold_WADDR6_WCLKS_posedge_posedge,
                             thold_WADDR6_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WCLKS_posedge,
                             TmDt_WADDR6_WCLKS_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR6_WCLKS_negedge_posedge,
                             tsetup_WADDR6_WCLKS_negedge_posedge,
                             thold_WADDR6_WCLKS_negedge_posedge,
                             thold_WADDR6_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WCLKS_posedge,
                             TmDt_WADDR7_WCLKS_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR7_WCLKS_posedge_posedge,
                             tsetup_WADDR7_WCLKS_posedge_posedge,
                             thold_WADDR7_WCLKS_posedge_posedge,
                             thold_WADDR7_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WCLKS_posedge,
                             TmDt_WADDR7_WCLKS_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR7_WCLKS_negedge_posedge,
                             tsetup_WADDR7_WCLKS_negedge_posedge,
                             thold_WADDR7_WCLKS_negedge_posedge,
                             thold_WADDR7_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_posedge_posedge,
                             tsetup_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_negedge_posedge,
                             tsetup_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_posedge_posedge,
                             tsetup_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_negedge_posedge,
                             tsetup_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_posedge_posedge,
                             tsetup_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_negedge_posedge,
                             tsetup_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_posedge_posedge,
                             tsetup_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_negedge_posedge,
                             tsetup_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_posedge_posedge,
                             tsetup_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_negedge_posedge,
                             tsetup_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_posedge_posedge,
                             tsetup_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_negedge_posedge,
                             tsetup_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_posedge_posedge,
                             tsetup_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_negedge_posedge,
                             tsetup_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_posedge_posedge,
                             tsetup_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_negedge_posedge,
                             tsetup_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_posedge_posedge,
                             tsetup_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_negedge_posedge,
                             tsetup_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

 -- setup hold WEN, WBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_posedge_posedge,
                             tsetup_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_negedge_posedge,
                             tsetup_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

  --   Period of WCLK
      VitalPeriodPulseCheck ( Pviol_WCLKS,
                              PeriodData_WCLKS,
                              WCLKS_ipd, "WCLKS",
                              0.0 ns,
                              tperiod_WCLKS,
                              tpw_WCLKS_posedge,
                              tpw_WCLKS_negedge,
                              (To_X01(WBLKB_ipd) = '0') AND (To_X01(WRB_ipd) = '0'),
                             InstancePath & "/RAM256x9SA",
                              True,
                              True,
                              WARNING
                              );
   ------------------------------------------------------------
   --        Timing Checking for Read and write conflict     --
   ------------------------------------------------------------
       VitalSetupHoldCheck ( Tviol_RDB_WCLKS_posedge,
                             TmDt_RDB_WCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_RDB_WCLKS_negedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBint) = '0') AND (To_X01(RBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_WCLKS_negedge,
                             TmDt_RDB_WCLKS_negedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RDB_WCLKS_posedge_negedge,
                             0.0 ns,
                             (To_X01(WBint) = '0') AND (To_X01(RBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_WCLKS_posedge,
                             TmDt_RBLKB_WCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_RBLKB_WCLKS_negedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBint) = '0') AND (To_X01(RDB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_WCLKS_negedge,
                             TmDt_RBLKB_WCLKS_negedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RBLKB_WCLKS_posedge_negedge,
                             0.0 ns,
                             (To_X01(WBint) = '0') AND (To_X01(RDB_ipd) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WCLKS_negedge,
                             TmDt_RADDR0_WCLKS_negedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR0_WCLKS_posedge_negedge,
                             thold_RADDR0_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WCLKS_posedge,
                             TmDt_RADDR0_WCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_WCLKS_posedge_posedge,
                             tsetup_RADDR0_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WCLKS_negedge,
                             TmDt_RADDR0_WCLKS_negedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR0_WCLKS_negedge_negedge,
                             thold_RADDR0_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WCLKS_posedge,
                             TmDt_RADDR0_WCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_WCLKS_negedge_posedge,
                             tsetup_RADDR0_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WCLKS_negedge,
                             TmDt_RADDR1_WCLKS_negedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR1_WCLKS_posedge_negedge,
                             thold_RADDR1_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WCLKS_posedge,
                             TmDt_RADDR1_WCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_WCLKS_posedge_posedge,
                             tsetup_RADDR1_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WCLKS_negedge,
                             TmDt_RADDR1_WCLKS_negedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR1_WCLKS_negedge_negedge,
                             thold_RADDR1_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WCLKS_posedge,
                             TmDt_RADDR1_WCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_WCLKS_negedge_posedge,
                             tsetup_RADDR1_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WCLKS_negedge,
                             TmDt_RADDR2_WCLKS_negedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR2_WCLKS_posedge_negedge,
                             thold_RADDR2_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WCLKS_posedge,
                             TmDt_RADDR2_WCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_WCLKS_posedge_posedge,
                             tsetup_RADDR2_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WCLKS_negedge,
                             TmDt_RADDR2_WCLKS_negedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR2_WCLKS_negedge_negedge,
                             thold_RADDR2_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WCLKS_posedge,
                             TmDt_RADDR2_WCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_WCLKS_negedge_posedge,
                             tsetup_RADDR2_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WCLKS_negedge,
                             TmDt_RADDR3_WCLKS_negedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR3_WCLKS_posedge_negedge,
                             thold_RADDR3_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WCLKS_posedge,
                             TmDt_RADDR3_WCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_WCLKS_posedge_posedge,
                             tsetup_RADDR3_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WCLKS_negedge,
                             TmDt_RADDR3_WCLKS_negedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR3_WCLKS_negedge_negedge,
                             thold_RADDR3_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WCLKS_posedge,
                             TmDt_RADDR3_WCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_WCLKS_negedge_posedge,
                             tsetup_RADDR3_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WCLKS_negedge,
                             TmDt_RADDR4_WCLKS_negedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR4_WCLKS_posedge_negedge,
                             thold_RADDR4_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WCLKS_posedge,
                             TmDt_RADDR4_WCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_WCLKS_posedge_posedge,
                             tsetup_RADDR4_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WCLKS_negedge,
                             TmDt_RADDR4_WCLKS_negedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR4_WCLKS_negedge_negedge,
                             thold_RADDR4_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WCLKS_posedge,
                             TmDt_RADDR4_WCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_WCLKS_negedge_posedge,
                             tsetup_RADDR4_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WCLKS_negedge,
                             TmDt_RADDR5_WCLKS_negedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR5_WCLKS_posedge_negedge,
                             thold_RADDR5_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WCLKS_posedge,
                             TmDt_RADDR5_WCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_WCLKS_posedge_posedge,
                             tsetup_RADDR5_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WCLKS_negedge,
                             TmDt_RADDR5_WCLKS_negedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR5_WCLKS_negedge_negedge,
                             thold_RADDR5_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WCLKS_posedge,
                             TmDt_RADDR5_WCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_WCLKS_negedge_posedge,
                             tsetup_RADDR5_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WCLKS_negedge,
                             TmDt_RADDR6_WCLKS_negedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR6_WCLKS_posedge_negedge,
                             thold_RADDR6_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WCLKS_posedge,
                             TmDt_RADDR6_WCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_WCLKS_posedge_posedge,
                             tsetup_RADDR6_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WCLKS_negedge,
                             TmDt_RADDR6_WCLKS_negedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR6_WCLKS_negedge_negedge,
                             thold_RADDR6_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WCLKS_posedge,
                             TmDt_RADDR6_WCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_WCLKS_negedge_posedge,
                             tsetup_RADDR6_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WCLKS_negedge,
                             TmDt_RADDR7_WCLKS_negedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR7_WCLKS_posedge_negedge,
                             thold_RADDR7_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WCLKS_posedge,
                             TmDt_RADDR7_WCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_WCLKS_posedge_posedge,
                             tsetup_RADDR7_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WCLKS_negedge,
                             TmDt_RADDR7_WCLKS_negedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR7_WCLKS_negedge_negedge,
                             thold_RADDR7_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WCLKS_posedge,
                             TmDt_RADDR7_WCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_WCLKS_negedge_posedge,
                             tsetup_RADDR7_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SA",
                             True,
                             True,
                             WARNING
                             );

 end if;

   ------------------------------------------------------------
   --    wpe output                                           -
   ------------------------------------------------------------

   if ( PARODD_ipd'EVENT ) then
     RPE_zd := not RPE_zd;
     WPE_zd := not WPE_zd;
   end if;

   ------------------------------------------------------------
   --         WPE checking  block                            -
   ------------------------------------------------------------

     if ( WCLKS_ipd'EVENT ) then
        tmp_par  := DI7_delayed XOR DI6_delayed XOR DI5_delayed XOR DI4_delayed XOR DI3_delayed XOR DI2_delayed XOR DI1_delayed XOR DI0_delayed;
        tmp_par2 := (tmp_par xor DI8_delayed);

      if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
          ( TO_X01 ( WCLKS_ipd  ) = 'X' ) or 
          ( TO_X01 ( DI8_ipd )    = 'X' ) or
          ( TO_X01 ( DI7_ipd )    = 'X' ) or
          ( TO_X01 ( DI6_ipd )    = 'X' ) or
          ( TO_X01 ( DI5_ipd )    = 'X' ) or
          ( TO_X01 ( DI4_ipd )    = 'X' ) or
          ( TO_X01 ( DI3_ipd )    = 'X' ) or
          ( TO_X01 ( DI2_ipd )    = 'X' ) or
          ( TO_X01 ( DI1_ipd )    = 'X' ) or
          ( TO_X01 ( DI0_ipd )    = 'X' )
         ) then
        wpe_var  :=  'X';
      elsif ( TO_X01 ( WCLKS_ipd ) = '1' ) then
        if ( tmp_par2 /= PARODD_ipd ) then
          wpe_var  :=  '1';
        else
          wpe_var  :=  '0';
        end if;
      end if;
      RAM_di_int(8) := DI8_ipd;
      WPE_zd := wpe_var;
     end if;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

    if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
    end if; 

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

  if (TO_X01(WCLKS_ipd)='X') then
   if (TO_X01(WCLKS_previous) /= 'X') then
    assert false
    report ": WCLK unknown"
    severity Warning;
    end if;
   elsif (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      case TO_X01(WBint_delayed) is
          when '1' =>
            null;
          when '0' =>
           if(WADDR < 0) then
            if ((TO_X01(WADDR0_delayed) = 'X') and (TO_X01(WADDR0_previous) /= 'X')) then
             assert false
             report ": WADDR0 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR1_delayed) = 'X') and (TO_X01(WADDR1_previous) /= 'X')) then
             assert false
             report ": WADDR1 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR2_delayed) = 'X') and (TO_X01(WADDR2_previous) /= 'X')) then
             assert false
             report ": WADDR2 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR3_delayed) = 'X') and (TO_X01(WADDR3_previous) /= 'X')) then
             assert false
             report ": WADDR3 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR4_delayed) = 'X') and (TO_X01(WADDR4_previous) /= 'X')) then
             assert false
             report ": WADDR4 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR5_delayed) = 'X') and (TO_X01(WADDR5_previous) /= 'X')) then
             assert false
             report ": WADDR5 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR6_delayed) = 'X') and (TO_X01(WADDR6_previous) /= 'X')) then
             assert false
             report ": WADDR6 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR7_delayed) = 'X') and (TO_X01(WADDR7_previous) /= 'X')) then
             assert false
             report ": WADDR7 unknown"
             severity Warning;
            end if;
           else 
             RAM_di_int(7 downto 0) := DI7_delayed & DI6_delayed & DI5_delayed & DI4_delayed & DI3_delayed & DI2_delayed & DI1_delayed & DI0_delayed;
             memory_array(WADDR)  := RAM_di_int;
           end if;

         when others =>
          if (TO_X01(WBint_previous) /= 'X') then
             assert false
             report ": WRB or WBLKB unknown"
             severity Warning;
           end if;
      end case;
    end if;


 -----------------------------------------------------------
 --  Read Functional Section                              --
 -----------------------------------------------------------



-- Asynchronous RAM Read, Enable signal controlled;
  if ( RBint'event or RADDR0_ipd'event or RADDR1_ipd'event or 
       RADDR2_ipd'event or RADDR3_ipd'event or RADDR4_ipd'event or 
       RADDR5_ipd'event or RADDR6_ipd'event or RADDR7_ipd'event or
       WCLKS_ipd'event ) then
    if ( TO_X01 ( RBint ) = 'X' ) then
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          RPE_zd :='X';
          if (TO_X01(RBint_previous) /= 'X') then
             assert false
             report ": RDB or RBLKB unknown"
             severity Warning;
          end if;
    elsif ( RADDR < 0 ) then
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          RPE_zd :='X';
          if(TO_X01(RADDR0_ipd) = 'X') and (TO_X01(RADDR0_previous) /= 'X') then
             assert false
             report ": RADDR0 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR1_ipd) = 'X') and (TO_X01(RADDR1_previous) /= 'X') then
             assert false
             report ": RADDR1 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR2_ipd) = 'X') and (TO_X01(RADDR2_previous) /= 'X') then
             assert false
             report ": RADDR2 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR3_ipd) = 'X') and (TO_X01(RADDR3_previous) /= 'X') then
             assert false
             report ": RADDR3 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR4_ipd) = 'X') and (TO_X01(RADDR4_previous) /= 'X') then
             assert false
             report ": RADDR4 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR5_ipd) = 'X') and (TO_X01(RADDR5_previous) /= 'X') then
             assert false
             report ": RADDR5 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR6_ipd) = 'X') and (TO_X01(RADDR6_previous) /= 'X') then
             assert false
             report ": RADDR6 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR7_ipd) = 'X') and (TO_X01(RADDR7_previous) /= 'X') then
             assert false
             report ": RADDR7 unknown"
             severity Warning;
          end if;
    elsif ( WADDR = RADDR ) then
        if (( RBint'event AND ( TO_X01 ( RBint ) = '0' ) AND ( TO_X01 ( WCLKS_ipd ) = '0' )) OR
            ( WCLKS_ipd'event AND ( TO_X01 ( WCLKS_ipd ) = '0' ) AND ( TO_X01 ( RBint ) = '0' )) OR
            ( RBint'event AND ( TO_X01 ( RBint ) = '1' ) AND ( TO_X01 ( WBint ) = '0' )) OR
            (( not (( TO_X01 ( WBint ) = '0' ) and ( TO_X01 ( WCLKS_ipd ) = '1' ))) AND 
             ( TO_X01 ( RBint ) = '0' ) AND 
             ( RADDR0_ipd'event or RADDR1_ipd'event or 
               RADDR2_ipd'event or RADDR3_ipd'event or RADDR4_ipd'event or 
               RADDR5_ipd'event or RADDR6_ipd'event or RADDR7_ipd'event ))
           ) then
             DO0_zd := memory_array(RADDR)(0);
             DO1_zd := memory_array(RADDR)(1);
             DO2_zd := memory_array(RADDR)(2);
             DO3_zd := memory_array(RADDR)(3);
             DO4_zd := memory_array(RADDR)(4);
             DO5_zd := memory_array(RADDR)(5);
             DO6_zd := memory_array(RADDR)(6);
             DO7_zd := memory_array(RADDR)(7);
             DO8_zd := memory_array(RADDR)(8);
             do_par := DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR 
                       DO3_zd XOR DO2_zd XOR DO1_zd XOR DO0_zd;
             if (do_par = 'X') then
               RPE_zd := 'X';
             elsif ( TO_X01 ( PARODD_ipd ) = 'X' ) then
               RPE_zd := 'X';
             else
               if (do_par /= PARODD_ipd) then
                 RPE_zd := '1';
               else
                 RPE_zd :=  '0';
               end if;
             end if;
        end if;
    else -- WADDR /= RADDR
        if ((( TO_X01 ( RBint ) = '0' ) AND
            ( RADDR0_ipd'event or RADDR1_ipd'event or RADDR2_ipd'event or 
              RADDR3_ipd'event or RADDR4_ipd'event or RADDR5_ipd'event or 
              RADDR6_ipd'event or RADDR7_ipd'event )) OR
           ( RBint'event AND ( TO_X01 ( RBint ) = '0' )) OR
           (( TO_X01 ( RBint ) = '0' ) AND
            ( RADDR0_ipd'event or RADDR1_ipd'event or RADDR2_ipd'event or 
              RADDR3_ipd'event or RADDR4_ipd'event or RADDR5_ipd'event or 
              RADDR6_ipd'event or RADDR7_ipd'event ))
          ) then
             DO0_zd := memory_array(RADDR)(0);
             DO1_zd := memory_array(RADDR)(1);
             DO2_zd := memory_array(RADDR)(2);
             DO3_zd := memory_array(RADDR)(3);
             DO4_zd := memory_array(RADDR)(4);
             DO5_zd := memory_array(RADDR)(5);
             DO6_zd := memory_array(RADDR)(6);
             DO7_zd := memory_array(RADDR)(7);
             DO8_zd := memory_array(RADDR)(8);
             
             do_par := DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR 
                       DO3_zd XOR DO2_zd XOR DO1_zd XOR DO0_zd;
             if (do_par = 'X') then
               RPE_zd := 'X';
             elsif ( TO_X01 ( PARODD_ipd ) = 'X' ) then
               RPE_zd := 'X';
             else
               if (do_par /= PARODD_ipd) then
                 RPE_zd := '1';
               else
                 RPE_zd :=  '0';
               end if;
             end if;
        end if;
    end if;  -- WADDR /= RADDR
  end if;




  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       WCLKS_previous  := WCLKS_ipd;
       RBint_previous  := RBint;
       WBint_previous  := WBint_delayed;
       WBint_delayed   := WBint;
       DI0_delayed     := DI0_ipd;
       DI1_delayed     := DI1_ipd;
       DI2_delayed     := DI2_ipd;
       DI3_delayed     := DI3_ipd;
       DI4_delayed     := DI4_ipd;
       DI5_delayed     := DI5_ipd;
       DI6_delayed     := DI6_ipd;
       DI7_delayed     := DI7_ipd;
       DI8_delayed     := DI8_ipd;
       RADDR0_previous := RADDR0_ipd;
       RADDR1_previous := RADDR1_ipd;
       RADDR2_previous := RADDR2_ipd;
       RADDR3_previous := RADDR3_ipd;
       RADDR4_previous := RADDR4_ipd;
       RADDR5_previous := RADDR5_ipd;
       RADDR6_previous := RADDR6_ipd;
       RADDR7_previous := RADDR7_ipd;
       WADDR0_previous := WADDR0_delayed;
       WADDR0_delayed  := WADDR0_ipd;
       WADDR1_previous := WADDR1_delayed;
       WADDR1_delayed  := WADDR1_ipd;
       WADDR2_previous := WADDR2_delayed;
       WADDR2_delayed  := WADDR2_ipd;
       WADDR3_previous := WADDR3_delayed;
       WADDR3_delayed  := WADDR3_ipd;
       WADDR4_previous := WADDR4_delayed;
       WADDR4_delayed  := WADDR4_ipd;
       WADDR5_previous := WADDR5_delayed;
       WADDR5_delayed  := WADDR5_ipd;
       WADDR6_previous := WADDR6_delayed;
       WADDR6_delayed  := WADDR6_ipd;
       WADDR7_previous := WADDR7_delayed;
       WADDR7_delayed  := WADDR7_ipd;
       PARODD_previous := PARODD_delayed; 
       PARODD_delayed  := PARODD_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
           OutSignal     => DOS,
           GlitchData    => DOS_GlitchData,
           OutSignalName => "DOS",
           OutTemp       => DOS_zd,
           Paths  =>  (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),
           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
             OutSignal     => WPE,
             GlitchData    => WPE_GlitchData,
             OutSignalName => "WPE",
             OutTemp       => WPE_zd,
             Paths =>   (0 => (WCLKS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_WCLKS_WPE), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO0), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO0), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO0), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO0), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO0), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO0), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO0), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO0), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO0), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO1), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO1), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO1), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO1), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO1), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO1), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO1), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO1), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO1), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO2), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO2), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO2), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO2), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO2), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO2), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO2), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO2), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO2), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO3), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO3), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO3), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO3), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO3), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO3), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO3), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO3), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO3), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO4), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO4), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO4), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO4), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO4), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO4), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO4), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO4), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO4), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO5), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO5), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO5), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO5), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO5), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO5), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO5), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO5), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO5), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO6), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO6), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO6), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO6), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO6), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO6), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO6), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO6), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO6), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO7), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO7), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO7), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO7), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO7), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO7), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO7), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO7), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO7), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO8), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO8), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO8), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO8), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO8), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO8), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO8), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO8), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO8), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => RPE,
           GlitchData    => RPE_GlitchData,
           OutSignalName => "RPE",
           OutTemp       => RPE_zd,

           Paths  =>   (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_RPE), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_RPE), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_RPE), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_RPE), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_RPE), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_RPE), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_RPE), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_RPE), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_RPE), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_RPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
LIBRARY STD;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

USE std.textio.all;
USE ieee.std_logic_textio.all;
LIBRARY a500k;
USE a500k.all;

entity RAM256x9SAP is 

   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR0_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR1_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR2_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR3_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR4_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR5_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR6_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RADDR7_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpw_RDB_posedge	        : VitalDelayType := 0.000 ns;
 	tpw_RDB_negedge	        : VitalDelayType := 0.000 ns;
 	tperiod_RDB	        : VitalDelayType := 0.000 ns;
 	tpw_RBLKB_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RBLKB_negedge	: VitalDelayType := 0.000 ns;
 	tperiod_RBLKB	        : VitalDelayType := 0.000 ns;
 	tpw_RADDR0_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR0_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR1_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR2_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR3_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR4_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR5_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR6_negedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_posedge	: VitalDelayType := 0.000 ns;
 	tpw_RADDR7_negedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tpw_WCLKS_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                           : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_RDB_WCLKS_negedge_posedge       : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_WCLKS_negedge_posedge       : VitalDelayType := 0.000 ns;
 	tsetup_RADDR0_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR0_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR1_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR2_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR3_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR4_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR5_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR6_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_WCLKS_negedge_posedge     : VitalDelayType := 0.000 ns;
	tsetup_RADDR7_WCLKS_posedge_posedge     : VitalDelayType := 0.000 ns;
 	thold_RDB_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RBLKB_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR0_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR1_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR2_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR3_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR4_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR5_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR6_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_WCLKS_negedge_negedge	: VitalDelayType := 0.000 ns;
        thold_RADDR7_WCLKS_posedge_negedge	: VitalDelayType := 0.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   WCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');

ATTRIBUTE VITAL_LEVEL0 OF RAM256x9SAP : entity IS True ;
END RAM256x9SAP;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of RAM256x9SAP is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal WADDR0_ipd : std_ulogic := 'X';
   signal WADDR1_ipd : std_ulogic := 'X';
   signal WADDR2_ipd : std_ulogic := 'X';
   signal WADDR3_ipd : std_ulogic := 'X';
   signal WADDR4_ipd : std_ulogic := 'X';
   signal WADDR5_ipd : std_ulogic := 'X';
   signal WADDR6_ipd : std_ulogic := 'X';
   signal WADDR7_ipd : std_ulogic := 'X';
   signal RADDR0_ipd : std_ulogic := 'X';
   signal RADDR1_ipd : std_ulogic := 'X';
   signal RADDR2_ipd : std_ulogic := 'X';
   signal RADDR3_ipd : std_ulogic := 'X';
   signal RADDR4_ipd : std_ulogic := 'X';
   signal RADDR5_ipd : std_ulogic := 'X';
   signal RADDR6_ipd : std_ulogic := 'X';
   signal RADDR7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal WCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

	-- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';
   signal INIT_MEM   : std_logic:= '0';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic:= 'X';
   signal par_f2     : std_logic:= 'X';

 begin  --  VITAL_ACT
   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (WADDR0_ipd, WADDR0, VitalExtendToFillDelay(tipd_WADDR0));
   VitalWireDelay (WADDR1_ipd, WADDR1, VitalExtendToFillDelay(tipd_WADDR1));
   VitalWireDelay (WADDR2_ipd, WADDR2, VitalExtendToFillDelay(tipd_WADDR2));
   VitalWireDelay (WADDR3_ipd, WADDR3, VitalExtendToFillDelay(tipd_WADDR3));
   VitalWireDelay (WADDR4_ipd, WADDR4, VitalExtendToFillDelay(tipd_WADDR4));
   VitalWireDelay (WADDR5_ipd, WADDR5, VitalExtendToFillDelay(tipd_WADDR5));
   VitalWireDelay (WADDR6_ipd, WADDR6, VitalExtendToFillDelay(tipd_WADDR6));
   VitalWireDelay (WADDR7_ipd, WADDR7, VitalExtendToFillDelay(tipd_WADDR7));
   VitalWireDelay (RADDR0_ipd, RADDR0, VitalExtendToFillDelay(tipd_RADDR0));
   VitalWireDelay (RADDR1_ipd, RADDR1, VitalExtendToFillDelay(tipd_RADDR1));
   VitalWireDelay (RADDR2_ipd, RADDR2, VitalExtendToFillDelay(tipd_RADDR2));
   VitalWireDelay (RADDR3_ipd, RADDR3, VitalExtendToFillDelay(tipd_RADDR3));
   VitalWireDelay (RADDR4_ipd, RADDR4, VitalExtendToFillDelay(tipd_RADDR4));
   VitalWireDelay (RADDR5_ipd, RADDR5, VitalExtendToFillDelay(tipd_RADDR5));
   VitalWireDelay (RADDR6_ipd, RADDR6, VitalExtendToFillDelay(tipd_RADDR6));
   VitalWireDelay (RADDR7_ipd, RADDR7, VitalExtendToFillDelay(tipd_RADDR7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (WCLKS_ipd, WCLKS, VitalExtendToFillDelay(tipd_WCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

---------------------------------------------------------------
--                  Behavior Section                         --
---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);


    PROCESS
    BEGIN
      INIT_MEM <= '1';
      WAIT;
    END PROCESS;

    VITALBehavior : process (INIT_MEM, 
                          RADDR0_ipd, RADDR1_ipd, RADDR2_ipd, RADDR3_ipd, RADDR4_ipd, RADDR5_ipd, RADDR6_ipd, RADDR7_ipd, 
                          WADDR0_ipd, WADDR1_ipd, WADDR2_ipd, WADDR3_ipd, WADDR4_ipd, WADDR5_ipd, WADDR6_ipd, WADDR7_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          WCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd 
                          )

    -- some internal veriable declaration
     variable RAM_di_int         : std_logic_vector(8 downto 0);
     variable memory_array       : MEM_TYPE := (others =>(others => 'X'));
     variable do_par             : std_logic:= 'X';
     variable tmp_par            : std_logic:= 'X';
     variable tmp_par2           : std_logic:= 'X';
     variable wpe_var            : std_logic:= 'X';

     --  Read Timing Check Results
     variable PeriodData_RDB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RDB                  : X01                 := '0';
     variable PeriodData_RBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RBLKB                : X01                  := '0';
     variable PeriodData_RADDR0          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR0               : X01                 := '0';
     variable PeriodData_RADDR1          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR1               : X01                 := '0';
     variable PeriodData_RADDR2          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR2               : X01                 := '0';
     variable PeriodData_RADDR3          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR3               : X01                 := '0';
     variable PeriodData_RADDR4          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR4               : X01                 := '0';
     variable PeriodData_RADDR5          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR5               : X01                 := '0';
     variable PeriodData_RADDR6          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR6               : X01                 := '0';
     variable PeriodData_RADDR7          : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RADDR7               : X01                 := '0';
     variable Tviol_WADDR0_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR0_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR1_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR2_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR3_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR4_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR5_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR6_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR7_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI0_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI1_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI2_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI3_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI4_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI5_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI6_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI7_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI8_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_WCLKS_posedge    : X01                 := '0';
     variable TmDt_WRB_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_WCLKS_posedge  : X01                 := '0';
     variable TmDt_WBLKB_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WCLKS                : X01                 := '0';
     variable Tviol_RDB_WCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_WCLKS_posedge    : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_WCLKS_negedge    : X01                 := '0';
     variable TmDt_RDB_WCLKS_negedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_WCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_WCLKS_negedge  : X01                 := '0';
     variable TmDt_RBLKB_WCLKS_negedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR0_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR0_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR0_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR0_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR1_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR1_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR2_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR2_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR3_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR3_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR4_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR4_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR5_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR5_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR6_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR6_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_WCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR7_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_WCLKS_negedge : X01                 := '0';
     variable TmDt_RADDR7_WCLKS_negedge  : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results

     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     variable DO0_zd : std_ulogic;
     variable DO1_zd : std_ulogic;
     variable DO2_zd : std_ulogic;
     variable DO3_zd : std_ulogic;
     variable DO4_zd : std_ulogic;
     variable DO5_zd : std_ulogic;
     variable DO6_zd : std_ulogic;
     variable DO7_zd : std_ulogic;
     variable DO8_zd : std_ulogic;
     variable RPE_zd : std_ulogic;
     variable WPE_zd : std_ulogic;
     variable DOS_zd : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData  : VitalGlitchDataType;
     variable DO1_GlitchData  : VitalGlitchDataType;
     variable DO2_GlitchData  : VitalGlitchDataType;
     variable DO3_GlitchData  : VitalGlitchDataType;
     variable DO4_GlitchData  : VitalGlitchDataType;
     variable DO5_GlitchData  : VitalGlitchDataType;
     variable DO6_GlitchData  : VitalGlitchDataType;
     variable DO7_GlitchData  : VitalGlitchDataType;
     variable DO8_GlitchData  : VitalGlitchDataType;
     variable DOS_GlitchData  : VitalGlitchDataType;

     -- last value variables
     variable WCLKS_previous  : std_ulogic := 'X';
     variable RBint_previous  : std_ulogic := 'X';
     variable WBint_delayed   : std_ulogic := 'X';
     variable WBint_previous  : std_ulogic := 'X';
     variable DIS_previous    : std_ulogic := 'X';
     variable DI0_delayed     : std_ulogic := 'X';
     variable DI1_delayed     : std_ulogic := 'X';
     variable DI2_delayed     : std_ulogic := 'X';
     variable DI3_delayed     : std_ulogic := 'X';
     variable DI4_delayed     : std_ulogic := 'X';
     variable DI5_delayed     : std_ulogic := 'X';
     variable DI6_delayed     : std_ulogic := 'X';
     variable DI7_delayed     : std_ulogic := 'X';
     variable DI8_delayed     : std_ulogic := 'X';
     variable RADDR0_previous : std_ulogic := 'X';
     variable RADDR1_previous : std_ulogic := 'X';
     variable RADDR2_previous : std_ulogic := 'X';
     variable RADDR3_previous : std_ulogic := 'X';
     variable RADDR4_previous : std_ulogic := 'X';
     variable RADDR5_previous : std_ulogic := 'X';
     variable RADDR6_previous : std_ulogic := 'X';
     variable RADDR7_previous : std_ulogic := 'X';
     variable WADDR0_delayed  : std_ulogic := 'X';
     variable WADDR1_delayed  : std_ulogic := 'X';
     variable WADDR2_delayed  : std_ulogic := 'X';
     variable WADDR3_delayed  : std_ulogic := 'X';
     variable WADDR4_delayed  : std_ulogic := 'X';
     variable WADDR5_delayed  : std_ulogic := 'X';
     variable WADDR6_delayed  : std_ulogic := 'X';
     variable WADDR7_delayed  : std_ulogic := 'X';
     variable WADDR0_previous : std_ulogic := 'X';
     variable WADDR1_previous : std_ulogic := 'X';
     variable WADDR2_previous : std_ulogic := 'X';
     variable WADDR3_previous : std_ulogic := 'X';
     variable WADDR4_previous : std_ulogic := 'X';
     variable WADDR5_previous : std_ulogic := 'X';
     variable WADDR6_previous : std_ulogic := 'X';
     variable WADDR7_previous : std_ulogic := 'X';

     variable PARODD_delayed  : std_ulogic := 'X';
     variable PARODD_previous : std_ulogic := 'X';
 
     variable inline    : LINE;
     variable indata    : std_logic_vector(8 downto 0);
     variable resdata   : std_logic_vector(8 downto 0);
     variable i         : integer:=0;
     file     memfile   : text;
     variable status         : file_open_status;
 
 begin -- process VITALBehavior

  -----------------------------------------------------------
  --    Initialize memory file from MEMORYFILE string      --
  -----------------------------------------------------------

  if ( INIT_MEM'EVENT and INIT_MEM = '1') then
    file_open(status, memfile, MEMORYFILE, read_mode);
    if ( status=open_ok ) then
      while((i < 256) and (not ENDFILE(memfile))) loop
        readline(memfile,inline);
        read(inline,indata);
        resdata := indata;
        memory_array(i) := resdata;
        i := i+1;
      end loop;
    else
      assert ( MEMORYFILE'length = 0 )
        report "Failed to open RAM256x9SAP memory initialization file in read mode"
        severity Note;
    end if;
    file_close(memfile);
  end if;


     if (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      WADDR := ((INT(WADDR7_delayed)*128)+(INT(WADDR6_delayed)*64)+(INT(
               WADDR5_delayed)*32) + (INT(WADDR4_delayed)*16) + 
               (INT(WADDR3_delayed)*8) + (INT(WADDR2_delayed)*4) + (INT(
               WADDR1_delayed)*2) + (INT(WADDR0_delayed)*1));
     end if;

   -- Convert Read Address Signal to Integer

      RADDR := ((INT(RADDR7_ipd)*128)+(INT(RADDR6_ipd)*64)+(INT(
               RADDR5_ipd)*32) + (INT(RADDR4_ipd)*16) + 
               (INT(RADDR3_ipd)*8) + (INT(RADDR2_ipd)*4) + (INT(
               RADDR1_ipd)*2) + (INT(RADDR0_ipd)*1));

if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

      VitalPeriodPulseCheck ( Pviol_RDB,
                              PeriodData_RDB,
                              RDB_ipd, "RDB",
                              0.0 ns,
                              tperiod_RDB,
                              tpw_RDB_posedge,
                              tpw_RDB_negedge,
                              (To_X01(RBLKB_ipd) = '0'),
                             InstancePath &"/RAM256x9SAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RBLKB,
                              PeriodData_RBLKB,
                              RBLKB_ipd, "RBLKB",
                              0.0 ns,
                              tperiod_RBLKB,
                              tpw_RBLKB_posedge,
                              tpw_RBLKB_negedge,
                              (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR0,
                              PeriodData_RADDR0,
                              RADDR0_ipd, "RADDR0",
                              0.0 ns,
                              tpw_RADDR0_posedge + tpw_RADDR0_posedge,
                              tpw_RADDR0_posedge,
                              tpw_RADDR0_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR1,
                              PeriodData_RADDR1,
                              RADDR1_ipd, "RADDR1",
                              0.0 ns,
                              tpw_RADDR1_posedge + tpw_RADDR1_posedge,
                              tpw_RADDR1_posedge,
                              tpw_RADDR1_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR2,
                              PeriodData_RADDR2,
                              RADDR2_ipd, "RADDR2",
                              0.0 ns,
                              tpw_RADDR2_posedge + tpw_RADDR2_posedge,
                              tpw_RADDR2_posedge,
                              tpw_RADDR2_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR3,
                              PeriodData_RADDR3,
                              RADDR3_ipd, "RADDR3",
                              0.0 ns,
                              tpw_RADDR3_posedge + tpw_RADDR3_posedge,
                              tpw_RADDR3_posedge,
                              tpw_RADDR3_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR4,
                              PeriodData_RADDR4,
                              RADDR4_ipd, "RADDR4",
                              0.0 ns,
                              tpw_RADDR4_posedge + tpw_RADDR4_posedge,
                              tpw_RADDR4_posedge,
                              tpw_RADDR4_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR5,
                              PeriodData_RADDR5,
                              RADDR5_ipd, "RADDR5",
                              0.0 ns,
                              tpw_RADDR5_posedge + tpw_RADDR5_posedge,
                              tpw_RADDR5_posedge,
                              tpw_RADDR5_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR6,
                              PeriodData_RADDR6,
                              RADDR6_ipd, "RADDR6",
                              0.0 ns,
                              tpw_RADDR6_posedge + tpw_RADDR6_posedge,
                              tpw_RADDR6_posedge,
                              tpw_RADDR6_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RADDR7,
                              PeriodData_RADDR7,
                              RADDR7_ipd, "RADDR7",
                              0.0 ns,
                              tpw_RADDR7_posedge + tpw_RADDR7_posedge,
                              tpw_RADDR7_posedge,
                              tpw_RADDR7_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SAP",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_WADDR0_WCLKS_posedge,
                             TmDt_WADDR0_WCLKS_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR0_WCLKS_posedge_posedge,
                             tsetup_WADDR0_WCLKS_posedge_posedge,
                             thold_WADDR0_WCLKS_posedge_posedge,
                             thold_WADDR0_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WCLKS_posedge,
                             TmDt_WADDR0_WCLKS_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR0_WCLKS_negedge_posedge,
                             tsetup_WADDR0_WCLKS_negedge_posedge,
                             thold_WADDR0_WCLKS_negedge_posedge,
                             thold_WADDR0_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WCLKS_posedge,
                             TmDt_WADDR1_WCLKS_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR1_WCLKS_posedge_posedge,
                             tsetup_WADDR1_WCLKS_posedge_posedge,
                             thold_WADDR1_WCLKS_posedge_posedge,
                             thold_WADDR1_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WCLKS_posedge,
                             TmDt_WADDR1_WCLKS_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR1_WCLKS_negedge_posedge,
                             tsetup_WADDR1_WCLKS_negedge_posedge,
                             thold_WADDR1_WCLKS_negedge_posedge,
                             thold_WADDR1_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WCLKS_posedge,
                             TmDt_WADDR2_WCLKS_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR2_WCLKS_posedge_posedge,
                             tsetup_WADDR2_WCLKS_posedge_posedge,
                             thold_WADDR2_WCLKS_posedge_posedge,
                             thold_WADDR2_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WCLKS_posedge,
                             TmDt_WADDR2_WCLKS_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR2_WCLKS_negedge_posedge,
                             tsetup_WADDR2_WCLKS_negedge_posedge,
                             thold_WADDR2_WCLKS_negedge_posedge,
                             thold_WADDR2_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WCLKS_posedge,
                             TmDt_WADDR3_WCLKS_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR3_WCLKS_posedge_posedge,
                             tsetup_WADDR3_WCLKS_posedge_posedge,
                             thold_WADDR3_WCLKS_posedge_posedge,
                             thold_WADDR3_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WCLKS_posedge,
                             TmDt_WADDR3_WCLKS_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR3_WCLKS_negedge_posedge,
                             tsetup_WADDR3_WCLKS_negedge_posedge,
                             thold_WADDR3_WCLKS_negedge_posedge,
                             thold_WADDR3_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WCLKS_posedge,
                             TmDt_WADDR4_WCLKS_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR4_WCLKS_posedge_posedge,
                             tsetup_WADDR4_WCLKS_posedge_posedge,
                             thold_WADDR4_WCLKS_posedge_posedge,
                             thold_WADDR4_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WCLKS_posedge,
                             TmDt_WADDR4_WCLKS_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR4_WCLKS_negedge_posedge,
                             tsetup_WADDR4_WCLKS_negedge_posedge,
                             thold_WADDR4_WCLKS_negedge_posedge,
                             thold_WADDR4_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WCLKS_posedge,
                             TmDt_WADDR5_WCLKS_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR5_WCLKS_posedge_posedge,
                             tsetup_WADDR5_WCLKS_posedge_posedge,
                             thold_WADDR5_WCLKS_posedge_posedge,
                             thold_WADDR5_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WCLKS_posedge,
                             TmDt_WADDR5_WCLKS_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR5_WCLKS_negedge_posedge,
                             tsetup_WADDR5_WCLKS_negedge_posedge,
                             thold_WADDR5_WCLKS_negedge_posedge,
                             thold_WADDR5_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WCLKS_posedge,
                             TmDt_WADDR6_WCLKS_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR6_WCLKS_posedge_posedge,
                             tsetup_WADDR6_WCLKS_posedge_posedge,
                             thold_WADDR6_WCLKS_posedge_posedge,
                             thold_WADDR6_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WCLKS_posedge,
                             TmDt_WADDR6_WCLKS_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR6_WCLKS_negedge_posedge,
                             tsetup_WADDR6_WCLKS_negedge_posedge,
                             thold_WADDR6_WCLKS_negedge_posedge,
                             thold_WADDR6_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WCLKS_posedge,
                             TmDt_WADDR7_WCLKS_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR7_WCLKS_posedge_posedge,
                             tsetup_WADDR7_WCLKS_posedge_posedge,
                             thold_WADDR7_WCLKS_posedge_posedge,
                             thold_WADDR7_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WCLKS_posedge,
                             TmDt_WADDR7_WCLKS_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR7_WCLKS_negedge_posedge,
                             tsetup_WADDR7_WCLKS_negedge_posedge,
                             thold_WADDR7_WCLKS_negedge_posedge,
                             thold_WADDR7_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_posedge_posedge,
                             tsetup_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_negedge_posedge,
                             tsetup_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_posedge_posedge,
                             tsetup_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_negedge_posedge,
                             tsetup_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_posedge_posedge,
                             tsetup_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_negedge_posedge,
                             tsetup_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_posedge_posedge,
                             tsetup_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_negedge_posedge,
                             tsetup_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_posedge_posedge,
                             tsetup_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_negedge_posedge,
                             tsetup_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_posedge_posedge,
                             tsetup_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_negedge_posedge,
                             tsetup_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_posedge_posedge,
                             tsetup_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_negedge_posedge,
                             tsetup_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_posedge_posedge,
                             tsetup_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_negedge_posedge,
                             tsetup_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_posedge_posedge,
                             tsetup_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_negedge_posedge,
                             tsetup_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

 -- setup hold WEN, WBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_posedge_posedge,
                             tsetup_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_negedge_posedge,
                             tsetup_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

  --   Period of WCLK
      VitalPeriodPulseCheck ( Pviol_WCLKS,
                              PeriodData_WCLKS,
                              WCLKS_ipd, "WCLKS",
                              0.0 ns,
                              tperiod_WCLKS,
                              tpw_WCLKS_posedge,
                              tpw_WCLKS_negedge,
                              (To_X01(WBLKB_ipd) = '0') AND (To_X01(WRB_ipd) = '0'),
                             InstancePath & "/RAM256x9SAP",
                              True,
                              True,
                              WARNING
                              );
   ------------------------------------------------------------
   --        Timing Checking for Read and write conflict     --
   ------------------------------------------------------------
       VitalSetupHoldCheck ( Tviol_RDB_WCLKS_posedge,
                             TmDt_RDB_WCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_RDB_WCLKS_negedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBint) = '0') AND (To_X01(RBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_WCLKS_negedge,
                             TmDt_RDB_WCLKS_negedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RDB_WCLKS_posedge_negedge,
                             0.0 ns,
                             (To_X01(WBint) = '0') AND (To_X01(RBLKB_ipd) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_WCLKS_posedge,
                             TmDt_RBLKB_WCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             tsetup_RBLKB_WCLKS_negedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             (To_X01(WBint) = '0') AND (To_X01(RDB_ipd) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_WCLKS_negedge,
                             TmDt_RBLKB_WCLKS_negedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RBLKB_WCLKS_posedge_negedge,
                             0.0 ns,
                             (To_X01(WBint) = '0') AND (To_X01(RDB_ipd) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WCLKS_negedge,
                             TmDt_RADDR0_WCLKS_negedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR0_WCLKS_posedge_negedge,
                             thold_RADDR0_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WCLKS_posedge,
                             TmDt_RADDR0_WCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_WCLKS_posedge_posedge,
                             tsetup_RADDR0_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WCLKS_negedge,
                             TmDt_RADDR0_WCLKS_negedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR0_WCLKS_negedge_negedge,
                             thold_RADDR0_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_WCLKS_posedge,
                             TmDt_RADDR0_WCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_WCLKS_negedge_posedge,
                             tsetup_RADDR0_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WCLKS_negedge,
                             TmDt_RADDR1_WCLKS_negedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR1_WCLKS_posedge_negedge,
                             thold_RADDR1_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WCLKS_posedge,
                             TmDt_RADDR1_WCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_WCLKS_posedge_posedge,
                             tsetup_RADDR1_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WCLKS_negedge,
                             TmDt_RADDR1_WCLKS_negedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR1_WCLKS_negedge_negedge,
                             thold_RADDR1_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_WCLKS_posedge,
                             TmDt_RADDR1_WCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_WCLKS_negedge_posedge,
                             tsetup_RADDR1_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WCLKS_negedge,
                             TmDt_RADDR2_WCLKS_negedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR2_WCLKS_posedge_negedge,
                             thold_RADDR2_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WCLKS_posedge,
                             TmDt_RADDR2_WCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_WCLKS_posedge_posedge,
                             tsetup_RADDR2_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WCLKS_negedge,
                             TmDt_RADDR2_WCLKS_negedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR2_WCLKS_negedge_negedge,
                             thold_RADDR2_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_WCLKS_posedge,
                             TmDt_RADDR2_WCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_WCLKS_negedge_posedge,
                             tsetup_RADDR2_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WCLKS_negedge,
                             TmDt_RADDR3_WCLKS_negedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR3_WCLKS_posedge_negedge,
                             thold_RADDR3_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WCLKS_posedge,
                             TmDt_RADDR3_WCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_WCLKS_posedge_posedge,
                             tsetup_RADDR3_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WCLKS_negedge,
                             TmDt_RADDR3_WCLKS_negedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR3_WCLKS_negedge_negedge,
                             thold_RADDR3_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_WCLKS_posedge,
                             TmDt_RADDR3_WCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_WCLKS_negedge_posedge,
                             tsetup_RADDR3_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WCLKS_negedge,
                             TmDt_RADDR4_WCLKS_negedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR4_WCLKS_posedge_negedge,
                             thold_RADDR4_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WCLKS_posedge,
                             TmDt_RADDR4_WCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_WCLKS_posedge_posedge,
                             tsetup_RADDR4_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WCLKS_negedge,
                             TmDt_RADDR4_WCLKS_negedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR4_WCLKS_negedge_negedge,
                             thold_RADDR4_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_WCLKS_posedge,
                             TmDt_RADDR4_WCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_WCLKS_negedge_posedge,
                             tsetup_RADDR4_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WCLKS_negedge,
                             TmDt_RADDR5_WCLKS_negedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR5_WCLKS_posedge_negedge,
                             thold_RADDR5_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WCLKS_posedge,
                             TmDt_RADDR5_WCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_WCLKS_posedge_posedge,
                             tsetup_RADDR5_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WCLKS_negedge,
                             TmDt_RADDR5_WCLKS_negedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR5_WCLKS_negedge_negedge,
                             thold_RADDR5_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_WCLKS_posedge,
                             TmDt_RADDR5_WCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_WCLKS_negedge_posedge,
                             tsetup_RADDR5_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WCLKS_negedge,
                             TmDt_RADDR6_WCLKS_negedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR6_WCLKS_posedge_negedge,
                             thold_RADDR6_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WCLKS_posedge,
                             TmDt_RADDR6_WCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_WCLKS_posedge_posedge,
                             tsetup_RADDR6_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WCLKS_negedge,
                             TmDt_RADDR6_WCLKS_negedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR6_WCLKS_negedge_negedge,
                             thold_RADDR6_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_WCLKS_posedge,
                             TmDt_RADDR6_WCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_WCLKS_negedge_posedge,
                             tsetup_RADDR6_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WCLKS_negedge,
                             TmDt_RADDR7_WCLKS_negedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR7_WCLKS_posedge_negedge,
                             thold_RADDR7_WCLKS_posedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WCLKS_posedge,
                             TmDt_RADDR7_WCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_WCLKS_posedge_posedge,
                             tsetup_RADDR7_WCLKS_posedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WCLKS_negedge,
                             TmDt_RADDR7_WCLKS_negedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             0.0 ns, 
                             0.0 ns, 
                             thold_RADDR7_WCLKS_negedge_negedge,
                             thold_RADDR7_WCLKS_negedge_negedge,
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '\',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_WCLKS_posedge,
                             TmDt_RADDR7_WCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_WCLKS_negedge_posedge,
                             tsetup_RADDR7_WCLKS_negedge_posedge,
                             0.0 ns, 
                             0.0 ns, 
                             (To_X01(WBint) = '0') AND (To_X01(RBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SAP",
                             True,
                             True,
                             WARNING
                             );

 end if;

   ------------------------------------------------------------
   --         WPE generating  block                            -
   ------------------------------------------------------------

     if ( WCLKS_ipd'EVENT ) then
        tmp_par  := DI7_delayed XOR DI6_delayed XOR DI5_delayed XOR DI4_delayed XOR DI3_delayed XOR DI2_delayed XOR DI1_delayed XOR DI0_delayed;
      if (( TO_X01 ( PARODD_ipd ) = 'X' ) or
          ( TO_X01 ( WCLKS_ipd  ) = 'X' ) or
          ( TO_X01 ( DI7_ipd )    = 'X' ) or
          ( TO_X01 ( DI6_ipd )    = 'X' ) or
          ( TO_X01 ( DI5_ipd )    = 'X' ) or
          ( TO_X01 ( DI4_ipd )    = 'X' ) or
          ( TO_X01 ( DI3_ipd )    = 'X' ) or
          ( TO_X01 ( DI2_ipd )    = 'X' ) or
          ( TO_X01 ( DI1_ipd )    = 'X' ) or
          ( TO_X01 ( DI0_ipd )    = 'X' )
         ) then
        wpe_var  :=  'X';
      elsif ( TO_X01 ( WCLKS_ipd ) = '1' ) then
        if ( tmp_par /= PARODD_ipd ) then
          wpe_var  :=  '1';
        else
          wpe_var  :=  '0';
        end if;
      end if;
        RAM_di_int(8) := wpe_var;
        WPE_zd := wpe_var;
     end if;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

    if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
    end if; 

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

  if (TO_X01(WCLKS_ipd)='X') then
   if (TO_X01(WCLKS_previous) /= 'X') then
    assert false
    report ": WCLK unknown"
    severity Warning;
    end if;
   elsif (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      case TO_X01(WBint_delayed) is
          when '1' =>
            null;
          when '0' =>
           if(WADDR < 0) then
            if ((TO_X01(WADDR0_delayed) = 'X') and (TO_X01(WADDR0_previous) /= 'X')) then
             assert false
             report ": WADDR0 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR1_delayed) = 'X') and (TO_X01(WADDR1_previous) /= 'X')) then
             assert false
             report ": WADDR1 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR2_delayed) = 'X') and (TO_X01(WADDR2_previous) /= 'X')) then
             assert false
             report ": WADDR2 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR3_delayed) = 'X') and (TO_X01(WADDR3_previous) /= 'X')) then
             assert false
             report ": WADDR3 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR4_delayed) = 'X') and (TO_X01(WADDR4_previous) /= 'X')) then
             assert false
             report ": WADDR4 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR5_delayed) = 'X') and (TO_X01(WADDR5_previous) /= 'X')) then
             assert false
             report ": WADDR5 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR6_delayed) = 'X') and (TO_X01(WADDR6_previous) /= 'X')) then
             assert false
             report ": WADDR6 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR7_delayed) = 'X') and (TO_X01(WADDR7_previous) /= 'X')) then
             assert false
             report ": WADDR7 unknown"
             severity Warning;
            end if;
           else 
             RAM_di_int(7 downto 0) := DI7_delayed & DI6_delayed & DI5_delayed & DI4_delayed & DI3_delayed & DI2_delayed & DI1_delayed & DI0_delayed;
             memory_array(WADDR)  := RAM_di_int;
           end if;

         when others =>
          if (TO_X01(WBint_previous) /= 'X') then
             assert false
             report ": WRB or WBLKB unknown"
             severity Warning;
           end if;
      end case;
    end if;


 -----------------------------------------------------------
 --  Read Functional Section                              --
 -----------------------------------------------------------



-- Asynchronous RAM Read, Enable signal controlled;

  if ( RBint'event or RADDR0_ipd'event or RADDR1_ipd'event or 
       RADDR2_ipd'event or RADDR3_ipd'event or RADDR4_ipd'event or 
       RADDR5_ipd'event or RADDR6_ipd'event or RADDR7_ipd'event or
       WCLKS_ipd'event ) then
    if ( TO_X01 ( RBint ) = 'X' ) then
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          if (TO_X01(RBint_previous) /= 'X') then
             assert false
             report ": RDB or RBLKB unknown"
             severity Warning;
          end if;
    elsif ( RADDR < 0 ) then
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          if(TO_X01(RADDR0_ipd) = 'X') and (TO_X01(RADDR0_previous) /= 'X') then
             assert false
             report ": RADDR0 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR1_ipd) = 'X') and (TO_X01(RADDR1_previous) /= 'X') then
             assert false
             report ": RADDR1 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR2_ipd) = 'X') and (TO_X01(RADDR2_previous) /= 'X') then
             assert false
             report ": RADDR2 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR3_ipd) = 'X') and (TO_X01(RADDR3_previous) /= 'X') then
             assert false
             report ": RADDR3 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR4_ipd) = 'X') and (TO_X01(RADDR4_previous) /= 'X') then
             assert false
             report ": RADDR4 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR5_ipd) = 'X') and (TO_X01(RADDR5_previous) /= 'X') then
             assert false
             report ": RADDR5 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR6_ipd) = 'X') and (TO_X01(RADDR6_previous) /= 'X') then
             assert false
             report ": RADDR6 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR7_ipd) = 'X') and (TO_X01(RADDR7_previous) /= 'X') then
             assert false
             report ": RADDR7 unknown"
             severity Warning;
          end if;
    elsif ( WADDR = RADDR ) then
        if (( RBint'event AND ( TO_X01 ( RBint ) = '0' ) AND ( TO_X01 ( WCLKS_ipd ) = '0' )) OR
            ( WCLKS_ipd'event AND ( TO_X01 ( WCLKS_ipd ) = '0' ) AND ( TO_X01 ( RBint ) = '0' )) OR
            ( RBint'event AND ( TO_X01 ( RBint ) = '1' ) AND ( TO_X01 ( WBint ) = '0' )) OR
            (( not (( TO_X01 ( WBint ) = '0' ) and ( TO_X01 ( WCLKS_ipd ) = '1' ))) AND 
             ( TO_X01 ( RBint ) = '0' ) AND 
             ( RADDR0_ipd'event or RADDR1_ipd'event or 
               RADDR2_ipd'event or RADDR3_ipd'event or RADDR4_ipd'event or 
               RADDR5_ipd'event or RADDR6_ipd'event or RADDR7_ipd'event ))
           ) then
             DO0_zd := memory_array(RADDR)(0);
             DO1_zd := memory_array(RADDR)(1);
             DO2_zd := memory_array(RADDR)(2);
             DO3_zd := memory_array(RADDR)(3);
             DO4_zd := memory_array(RADDR)(4);
             DO5_zd := memory_array(RADDR)(5);
             DO6_zd := memory_array(RADDR)(6);
             DO7_zd := memory_array(RADDR)(7);
             DO8_zd := memory_array(RADDR)(8);
             do_par := DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR 
                       DO3_zd XOR DO2_zd XOR DO1_zd XOR DO0_zd;
        end if;
    else -- WADDR /= RADDR
        if ((( TO_X01 ( RBint ) = '0' ) AND
            ( RADDR0_ipd'event or RADDR1_ipd'event or RADDR2_ipd'event or 
              RADDR3_ipd'event or RADDR4_ipd'event or RADDR5_ipd'event or 
              RADDR6_ipd'event or RADDR7_ipd'event )) OR
           ( RBint'event AND ( TO_X01 ( RBint ) = '0' )) OR
           (( TO_X01 ( RBint ) = '0' ) AND
            ( RADDR0_ipd'event or RADDR1_ipd'event or RADDR2_ipd'event or 
              RADDR3_ipd'event or RADDR4_ipd'event or RADDR5_ipd'event or 
              RADDR6_ipd'event or RADDR7_ipd'event ))
          ) then
             DO0_zd := memory_array(RADDR)(0);
             DO1_zd := memory_array(RADDR)(1);
             DO2_zd := memory_array(RADDR)(2);
             DO3_zd := memory_array(RADDR)(3);
             DO4_zd := memory_array(RADDR)(4);
             DO5_zd := memory_array(RADDR)(5);
             DO6_zd := memory_array(RADDR)(6);
             DO7_zd := memory_array(RADDR)(7);
             DO8_zd := memory_array(RADDR)(8);
             
        end if;
    end if;  -- WADDR /= RADDR
  end if;


  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       WCLKS_previous  := WCLKS_ipd;
       RBint_previous  := RBint;
       WBint_previous  := WBint_delayed;
       WBint_delayed   := WBint;
       DI0_delayed     := DI0_ipd;
       DI1_delayed     := DI1_ipd;
       DI2_delayed     := DI2_ipd;
       DI3_delayed     := DI3_ipd;
       DI4_delayed     := DI4_ipd;
       DI5_delayed     := DI5_ipd;
       DI6_delayed     := DI6_ipd;
       DI7_delayed     := DI7_ipd;
       DI8_delayed     := DI8_ipd;
       RADDR0_previous := RADDR0_ipd;
       RADDR1_previous := RADDR1_ipd;
       RADDR2_previous := RADDR2_ipd;
       RADDR3_previous := RADDR3_ipd;
       RADDR4_previous := RADDR4_ipd;
       RADDR5_previous := RADDR5_ipd;
       RADDR6_previous := RADDR6_ipd;
       RADDR7_previous := RADDR7_ipd;
       WADDR0_previous := WADDR0_delayed;
       WADDR0_delayed  := WADDR0_ipd;
       WADDR1_previous := WADDR1_delayed;
       WADDR1_delayed  := WADDR1_ipd;
       WADDR2_previous := WADDR2_delayed;
       WADDR2_delayed  := WADDR2_ipd;
       WADDR3_previous := WADDR3_delayed;
       WADDR3_delayed  := WADDR3_ipd;
       WADDR4_previous := WADDR4_delayed;
       WADDR4_delayed  := WADDR4_ipd;
       WADDR5_previous := WADDR5_delayed;
       WADDR5_delayed  := WADDR5_ipd;
       WADDR6_previous := WADDR6_delayed;
       WADDR6_delayed  := WADDR6_ipd;
       WADDR7_previous := WADDR7_delayed;
       WADDR7_delayed  := WADDR7_ipd;
       PARODD_previous := PARODD_delayed; 
       PARODD_delayed  := PARODD_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
           OutSignal     => DOS,
           GlitchData    => DOS_GlitchData,
           OutSignalName => "DOS",
           OutTemp       => DOS_zd,
           Paths  =>  (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),
           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO0), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO0), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO0), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO0), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO0), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO0), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO0), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO0), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO0), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO1), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO1), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO1), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO1), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO1), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO1), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO1), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO1), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO1), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO2), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO2), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO2), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO2), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO2), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO2), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO2), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO2), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO2), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO3), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO3), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO3), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO3), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO3), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO3), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO3), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO3), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO3), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO4), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO4), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO4), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO4), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO4), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO4), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO4), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO4), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO4), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO5), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO5), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO5), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO5), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO5), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO5), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO5), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO5), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO5), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO6), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO6), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO6), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO6), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO6), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO6), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO6), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO6), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO6), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO7), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO7), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO7), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO7), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO7), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO7), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO7), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO7), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO7), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths  =>    (0 => (RADDR0_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR0_DO8), true),
                         1 => (RADDR1_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR1_DO8), true),
                         2 => (RADDR2_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR2_DO8), true),
                         3 => (RADDR3_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR3_DO8), true),
                         4 => (RADDR4_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR4_DO8), true),
                         5 => (RADDR5_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR5_DO8), true),
                         6 => (RADDR6_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR6_DO8), true),
                         7 => (RADDR7_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RADDR7_DO8), true),
                         8 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO8), true),
                         9 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
LIBRARY STD;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

USE std.textio.all;
USE ieee.std_logic_textio.all;
LIBRARY a500k;
USE a500k.all;

entity RAM256x9SST is 

   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_WCLKS_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tpw_WCLKS_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                           : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 7.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';
   WPE    :  OUT STD_LOGIC := 'X';
   RPE    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   WCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');

ATTRIBUTE VITAL_LEVEL0 OF RAM256x9SST : entity IS True ;
END RAM256x9SST;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of RAM256x9SST is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal WADDR0_ipd : std_ulogic := 'X';
   signal WADDR1_ipd : std_ulogic := 'X';
   signal WADDR2_ipd : std_ulogic := 'X';
   signal WADDR3_ipd : std_ulogic := 'X';
   signal WADDR4_ipd : std_ulogic := 'X';
   signal WADDR5_ipd : std_ulogic := 'X';
   signal WADDR6_ipd : std_ulogic := 'X';
   signal WADDR7_ipd : std_ulogic := 'X';
   signal RADDR0_ipd : std_ulogic := 'X';
   signal RADDR1_ipd : std_ulogic := 'X';
   signal RADDR2_ipd : std_ulogic := 'X';
   signal RADDR3_ipd : std_ulogic := 'X';
   signal RADDR4_ipd : std_ulogic := 'X';
   signal RADDR5_ipd : std_ulogic := 'X';
   signal RADDR6_ipd : std_ulogic := 'X';
   signal RADDR7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal WCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

	-- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';
   signal INIT_MEM   : std_logic:= '0';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic:= 'X';
   signal par_f2     : std_logic:= 'X';

 begin  --  VITAL_ACT
   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (WADDR0_ipd, WADDR0, VitalExtendToFillDelay(tipd_WADDR0));
   VitalWireDelay (WADDR1_ipd, WADDR1, VitalExtendToFillDelay(tipd_WADDR1));
   VitalWireDelay (WADDR2_ipd, WADDR2, VitalExtendToFillDelay(tipd_WADDR2));
   VitalWireDelay (WADDR3_ipd, WADDR3, VitalExtendToFillDelay(tipd_WADDR3));
   VitalWireDelay (WADDR4_ipd, WADDR4, VitalExtendToFillDelay(tipd_WADDR4));
   VitalWireDelay (WADDR5_ipd, WADDR5, VitalExtendToFillDelay(tipd_WADDR5));
   VitalWireDelay (WADDR6_ipd, WADDR6, VitalExtendToFillDelay(tipd_WADDR6));
   VitalWireDelay (WADDR7_ipd, WADDR7, VitalExtendToFillDelay(tipd_WADDR7));
   VitalWireDelay (RADDR0_ipd, RADDR0, VitalExtendToFillDelay(tipd_RADDR0));
   VitalWireDelay (RADDR1_ipd, RADDR1, VitalExtendToFillDelay(tipd_RADDR1));
   VitalWireDelay (RADDR2_ipd, RADDR2, VitalExtendToFillDelay(tipd_RADDR2));
   VitalWireDelay (RADDR3_ipd, RADDR3, VitalExtendToFillDelay(tipd_RADDR3));
   VitalWireDelay (RADDR4_ipd, RADDR4, VitalExtendToFillDelay(tipd_RADDR4));
   VitalWireDelay (RADDR5_ipd, RADDR5, VitalExtendToFillDelay(tipd_RADDR5));
   VitalWireDelay (RADDR6_ipd, RADDR6, VitalExtendToFillDelay(tipd_RADDR6));
   VitalWireDelay (RADDR7_ipd, RADDR7, VitalExtendToFillDelay(tipd_RADDR7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (WCLKS_ipd, WCLKS, VitalExtendToFillDelay(tipd_WCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

---------------------------------------------------------------
--                  Behavior Section                         --
---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);


    PROCESS
    BEGIN
      INIT_MEM <= '1';
      WAIT;
    END PROCESS;

    VITALBehavior : process (INIT_MEM, 
                          RADDR0_ipd, RADDR1_ipd, RADDR2_ipd, RADDR3_ipd, RADDR4_ipd, RADDR5_ipd, RADDR6_ipd, RADDR7_ipd, 
                          WADDR0_ipd, WADDR1_ipd, WADDR2_ipd, WADDR3_ipd, WADDR4_ipd, WADDR5_ipd, WADDR6_ipd, WADDR7_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd 
                          )

    -- some internal veriable declaration
     variable RAM_di_int         : std_logic_vector(8 downto 0);
     variable memory_array       : MEM_TYPE := (others =>(others => 'X'));
     variable do_par             : std_logic:= 'X';
     variable tmp_par            : std_logic:= 'X';
     variable tmp_par2           : std_logic:= 'X';
     variable wpe_var            : std_logic:= 'X';

     --  Read Timing Check Results
     variable Tviol_RADDR0_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR0_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR1_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR2_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR3_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR4_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR5_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR6_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR7_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable Tviol_WADDR0_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR0_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR1_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR2_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR3_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR4_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR5_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR6_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR7_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI0_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI1_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI2_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI3_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI4_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI5_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI6_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI7_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI8_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_WCLKS_posedge    : X01                 := '0';
     variable TmDt_WRB_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_WCLKS_posedge  : X01                 := '0';
     variable TmDt_WBLKB_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WCLKS                : X01                 := '0';
     variable Tviol_WCLKS_RCLKS_posedge  : X01                 := '0';
     variable TmDt_WCLKS_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results

     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     variable DO0_zd : std_ulogic;
     variable DO1_zd : std_ulogic;
     variable DO2_zd : std_ulogic;
     variable DO3_zd : std_ulogic;
     variable DO4_zd : std_ulogic;
     variable DO5_zd : std_ulogic;
     variable DO6_zd : std_ulogic;
     variable DO7_zd : std_ulogic;
     variable DO8_zd : std_ulogic;
     variable RPE_zd : std_ulogic;
     variable WPE_zd : std_ulogic;
     variable DOS_zd : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData  : VitalGlitchDataType;
     variable DO1_GlitchData  : VitalGlitchDataType;
     variable DO2_GlitchData  : VitalGlitchDataType;
     variable DO3_GlitchData  : VitalGlitchDataType;
     variable DO4_GlitchData  : VitalGlitchDataType;
     variable DO5_GlitchData  : VitalGlitchDataType;
     variable DO6_GlitchData  : VitalGlitchDataType;
     variable DO7_GlitchData  : VitalGlitchDataType;
     variable DO8_GlitchData  : VitalGlitchDataType;
     variable RPE_GlitchData  : VitalGlitchDataType;
     variable WPE_GlitchData  : VitalGlitchDataType;
     variable DOS_GlitchData  : VitalGlitchDataType;

     -- last value variables
     variable WCLKS_previous  : std_ulogic := 'X';
     variable RCLKS_previous  : std_ulogic := 'X';
     variable RBint_delayed   : std_ulogic := 'X';
     variable RBint_previous  : std_ulogic := 'X';
     variable WBint_delayed   : std_ulogic := 'X';
     variable WBint_previous  : std_ulogic := 'X';
     variable DIS_previous    : std_ulogic := 'X';
     variable DI0_delayed     : std_ulogic := 'X';
     variable DI1_delayed     : std_ulogic := 'X';
     variable DI2_delayed     : std_ulogic := 'X';
     variable DI3_delayed     : std_ulogic := 'X';
     variable DI4_delayed     : std_ulogic := 'X';
     variable DI5_delayed     : std_ulogic := 'X';
     variable DI6_delayed     : std_ulogic := 'X';
     variable DI7_delayed     : std_ulogic := 'X';
     variable DI8_delayed     : std_ulogic := 'X';
     variable RADDR0_delayed  : std_ulogic := 'X';
     variable RADDR1_delayed  : std_ulogic := 'X';
     variable RADDR2_delayed  : std_ulogic := 'X';
     variable RADDR3_delayed  : std_ulogic := 'X';
     variable RADDR4_delayed  : std_ulogic := 'X';
     variable RADDR5_delayed  : std_ulogic := 'X';
     variable RADDR6_delayed  : std_ulogic := 'X';
     variable RADDR7_delayed  : std_ulogic := 'X';
     variable RADDR0_previous : std_ulogic := 'X';
     variable RADDR1_previous : std_ulogic := 'X';
     variable RADDR2_previous : std_ulogic := 'X';
     variable RADDR3_previous : std_ulogic := 'X';
     variable RADDR4_previous : std_ulogic := 'X';
     variable RADDR5_previous : std_ulogic := 'X';
     variable RADDR6_previous : std_ulogic := 'X';
     variable RADDR7_previous : std_ulogic := 'X';
     variable WADDR0_delayed  : std_ulogic := 'X';
     variable WADDR1_delayed  : std_ulogic := 'X';
     variable WADDR2_delayed  : std_ulogic := 'X';
     variable WADDR3_delayed  : std_ulogic := 'X';
     variable WADDR4_delayed  : std_ulogic := 'X';
     variable WADDR5_delayed  : std_ulogic := 'X';
     variable WADDR6_delayed  : std_ulogic := 'X';
     variable WADDR7_delayed  : std_ulogic := 'X';
     variable WADDR0_previous : std_ulogic := 'X';
     variable WADDR1_previous : std_ulogic := 'X';
     variable WADDR2_previous : std_ulogic := 'X';
     variable WADDR3_previous : std_ulogic := 'X';
     variable WADDR4_previous : std_ulogic := 'X';
     variable WADDR5_previous : std_ulogic := 'X';
     variable WADDR6_previous : std_ulogic := 'X';
     variable WADDR7_previous : std_ulogic := 'X';

     variable PARODD_delayed  : std_ulogic := 'X';
     variable PARODD_previous : std_ulogic := 'X';

     variable inline    : LINE;
     variable indata    : std_logic_vector(8 downto 0);
     variable resdata   : std_logic_vector(8 downto 0);
     variable i         : integer:=0;
     file     memfile   : text;
     variable status         : file_open_status;

 begin -- process VITALBehavior


  -----------------------------------------------------------
  --    Initialize memory file from MEMORYFILE string      --
  -----------------------------------------------------------


  if ( INIT_MEM'EVENT and INIT_MEM = '1') then
    file_open(status, memfile, MEMORYFILE, read_mode);
    if ( status=open_ok ) then
      while((i < 256) and (not ENDFILE(memfile))) loop
        readline(memfile,inline);
        read(inline,indata);
        resdata := indata;
        memory_array(i) := resdata;
        i := i+1;
      end loop;
    else
      assert ( MEMORYFILE'length = 0 )
        report "Failed to open RAM256x9SST memory initialization file in read mode"
        severity Note;
    end if;
    file_close(memfile);
  end if;

     if (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      WADDR := ((INT(WADDR7_delayed)*128)+(INT(WADDR6_delayed)*64)+(INT(
               WADDR5_delayed)*32) + (INT(WADDR4_delayed)*16) + 
               (INT(WADDR3_delayed)*8) + (INT(WADDR2_delayed)*4) + (INT(
               WADDR1_delayed)*2) + (INT(WADDR0_delayed)*1));
     end if;

   -- Convert Read Address Signal to Integer
     if (RCLKS_ipd'EVENT AND RCLKS_ipd = '1') then
      RADDR := ((INT(RADDR7_delayed)*128)+(INT(RADDR6_delayed)*64)+(INT(
               RADDR5_delayed)*32) + (INT(RADDR4_delayed)*16) + 
               (INT(RADDR3_delayed)*8) + (INT(RADDR2_delayed)*4) + (INT(
               RADDR1_delayed)*2) + (INT(RADDR0_delayed)*1));
     end if;

if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

 -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SST",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_WADDR0_WCLKS_posedge,
                             TmDt_WADDR0_WCLKS_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR0_WCLKS_posedge_posedge,
                             tsetup_WADDR0_WCLKS_posedge_posedge,
                             thold_WADDR0_WCLKS_posedge_posedge,
                             thold_WADDR0_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WCLKS_posedge,
                             TmDt_WADDR0_WCLKS_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR0_WCLKS_negedge_posedge,
                             tsetup_WADDR0_WCLKS_negedge_posedge,
                             thold_WADDR0_WCLKS_negedge_posedge,
                             thold_WADDR0_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WCLKS_posedge,
                             TmDt_WADDR1_WCLKS_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR1_WCLKS_posedge_posedge,
                             tsetup_WADDR1_WCLKS_posedge_posedge,
                             thold_WADDR1_WCLKS_posedge_posedge,
                             thold_WADDR1_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WCLKS_posedge,
                             TmDt_WADDR1_WCLKS_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR1_WCLKS_negedge_posedge,
                             tsetup_WADDR1_WCLKS_negedge_posedge,
                             thold_WADDR1_WCLKS_negedge_posedge,
                             thold_WADDR1_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WCLKS_posedge,
                             TmDt_WADDR2_WCLKS_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR2_WCLKS_posedge_posedge,
                             tsetup_WADDR2_WCLKS_posedge_posedge,
                             thold_WADDR2_WCLKS_posedge_posedge,
                             thold_WADDR2_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WCLKS_posedge,
                             TmDt_WADDR2_WCLKS_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR2_WCLKS_negedge_posedge,
                             tsetup_WADDR2_WCLKS_negedge_posedge,
                             thold_WADDR2_WCLKS_negedge_posedge,
                             thold_WADDR2_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WCLKS_posedge,
                             TmDt_WADDR3_WCLKS_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR3_WCLKS_posedge_posedge,
                             tsetup_WADDR3_WCLKS_posedge_posedge,
                             thold_WADDR3_WCLKS_posedge_posedge,
                             thold_WADDR3_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WCLKS_posedge,
                             TmDt_WADDR3_WCLKS_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR3_WCLKS_negedge_posedge,
                             tsetup_WADDR3_WCLKS_negedge_posedge,
                             thold_WADDR3_WCLKS_negedge_posedge,
                             thold_WADDR3_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WCLKS_posedge,
                             TmDt_WADDR4_WCLKS_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR4_WCLKS_posedge_posedge,
                             tsetup_WADDR4_WCLKS_posedge_posedge,
                             thold_WADDR4_WCLKS_posedge_posedge,
                             thold_WADDR4_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WCLKS_posedge,
                             TmDt_WADDR4_WCLKS_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR4_WCLKS_negedge_posedge,
                             tsetup_WADDR4_WCLKS_negedge_posedge,
                             thold_WADDR4_WCLKS_negedge_posedge,
                             thold_WADDR4_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WCLKS_posedge,
                             TmDt_WADDR5_WCLKS_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR5_WCLKS_posedge_posedge,
                             tsetup_WADDR5_WCLKS_posedge_posedge,
                             thold_WADDR5_WCLKS_posedge_posedge,
                             thold_WADDR5_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WCLKS_posedge,
                             TmDt_WADDR5_WCLKS_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR5_WCLKS_negedge_posedge,
                             tsetup_WADDR5_WCLKS_negedge_posedge,
                             thold_WADDR5_WCLKS_negedge_posedge,
                             thold_WADDR5_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WCLKS_posedge,
                             TmDt_WADDR6_WCLKS_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR6_WCLKS_posedge_posedge,
                             tsetup_WADDR6_WCLKS_posedge_posedge,
                             thold_WADDR6_WCLKS_posedge_posedge,
                             thold_WADDR6_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WCLKS_posedge,
                             TmDt_WADDR6_WCLKS_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR6_WCLKS_negedge_posedge,
                             tsetup_WADDR6_WCLKS_negedge_posedge,
                             thold_WADDR6_WCLKS_negedge_posedge,
                             thold_WADDR6_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WCLKS_posedge,
                             TmDt_WADDR7_WCLKS_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR7_WCLKS_posedge_posedge,
                             tsetup_WADDR7_WCLKS_posedge_posedge,
                             thold_WADDR7_WCLKS_posedge_posedge,
                             thold_WADDR7_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WCLKS_posedge,
                             TmDt_WADDR7_WCLKS_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR7_WCLKS_negedge_posedge,
                             tsetup_WADDR7_WCLKS_negedge_posedge,
                             thold_WADDR7_WCLKS_negedge_posedge,
                             thold_WADDR7_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_posedge_posedge,
                             tsetup_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_negedge_posedge,
                             tsetup_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_posedge_posedge,
                             tsetup_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_negedge_posedge,
                             tsetup_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_posedge_posedge,
                             tsetup_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_negedge_posedge,
                             tsetup_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_posedge_posedge,
                             tsetup_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_negedge_posedge,
                             tsetup_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_posedge_posedge,
                             tsetup_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_negedge_posedge,
                             tsetup_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_posedge_posedge,
                             tsetup_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_negedge_posedge,
                             tsetup_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_posedge_posedge,
                             tsetup_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_negedge_posedge,
                             tsetup_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_posedge_posedge,
                             tsetup_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_negedge_posedge,
                             tsetup_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_posedge_posedge,
                             tsetup_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_negedge_posedge,
                             tsetup_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

 -- setup hold WEN, WBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_posedge_posedge,
                             tsetup_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_negedge_posedge,
                             tsetup_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

  --   Period of WCLK
      VitalPeriodPulseCheck ( Pviol_WCLKS,
                              PeriodData_WCLKS,
                              WCLKS_ipd, "WCLKS",
                              0.0 ns,
                              tperiod_WCLKS,
                              tpw_WCLKS_posedge,
                              tpw_WCLKS_negedge,
                              (To_X01(WBLKB_ipd) = '0') AND (To_X01(WRB_ipd) = '0'),
                             InstancePath & "/RAM256x9SST",
                              True,
                              True,
                              WARNING
                              );
   ------------------------------------------------------------
   --        Timing Checking for Read and write conflict     --
   ------------------------------------------------------------
       VitalSetupHoldCheck ( Tviol_WCLKS_RCLKS_posedge,
                             TmDt_WCLKS_RCLKS_posedge,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_WCLKS_RCLKS_posedge_posedge,
                             0.0 ns,
                             thold_WCLKS_RCLKS_posedge_posedge,
                             0.0 ns,
                             (To_X01(RBint) = '0') AND (To_X01(WBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SST",
                             True,
                             True,
                             WARNING
                             );

 end if;

   ------------------------------------------------------------
   --    wpe output                                           -
   ------------------------------------------------------------

   if ( PARODD_ipd'EVENT ) then
     RPE_zd := not RPE_zd;
     WPE_zd := not WPE_zd;
   end if;

   ------------------------------------------------------------
   --         WPE checking  block                            -
   ------------------------------------------------------------

     if ( WCLKS_ipd'EVENT ) then
        tmp_par  := DI7_delayed XOR DI6_delayed XOR DI5_delayed XOR DI4_delayed XOR DI3_delayed XOR DI2_delayed XOR DI1_delayed XOR DI0_delayed;
        tmp_par2 := (tmp_par xor DI8_delayed);

      if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
          ( TO_X01 ( WCLKS_ipd  ) = 'X' ) or 
          ( TO_X01 ( DI8_ipd )    = 'X' ) or
          ( TO_X01 ( DI7_ipd )    = 'X' ) or
          ( TO_X01 ( DI6_ipd )    = 'X' ) or
          ( TO_X01 ( DI5_ipd )    = 'X' ) or
          ( TO_X01 ( DI4_ipd )    = 'X' ) or
          ( TO_X01 ( DI3_ipd )    = 'X' ) or
          ( TO_X01 ( DI2_ipd )    = 'X' ) or
          ( TO_X01 ( DI1_ipd )    = 'X' ) or
          ( TO_X01 ( DI0_ipd )    = 'X' )
         ) then
        wpe_var  :=  'X';
      elsif ( TO_X01 ( WCLKS_ipd ) = '1' ) then
        if ( tmp_par2 /= PARODD_ipd ) then
          wpe_var  :=  '1';
        else
          wpe_var  :=  '0';
        end if;
      end if;
      RAM_di_int(8) := DI8_delayed;
      WPE_zd := wpe_var;
     end if;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

    if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
    end if; 

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

  if (TO_X01(WCLKS_ipd)='X') then
   if (TO_X01(WCLKS_previous) /= 'X') then
    assert false
    report ": WCLK unknown"
    severity Warning;
    end if;
   elsif (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      case TO_X01(WBint_delayed) is
          when '1' =>
            null;
          when '0' =>
           if(WADDR < 0) then
            if ((TO_X01(WADDR0_delayed) = 'X') and (TO_X01(WADDR0_previous) /= 'X')) then
             assert false
             report ": WADDR0 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR1_delayed) = 'X') and (TO_X01(WADDR1_previous) /= 'X')) then
             assert false
             report ": WADDR1 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR2_delayed) = 'X') and (TO_X01(WADDR2_previous) /= 'X')) then
             assert false
             report ": WADDR2 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR3_delayed) = 'X') and (TO_X01(WADDR3_previous) /= 'X')) then
             assert false
             report ": WADDR3 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR4_delayed) = 'X') and (TO_X01(WADDR4_previous) /= 'X')) then
             assert false
             report ": WADDR4 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR5_delayed) = 'X') and (TO_X01(WADDR5_previous) /= 'X')) then
             assert false
             report ": WADDR5 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR6_delayed) = 'X') and (TO_X01(WADDR6_previous) /= 'X')) then
             assert false
             report ": WADDR6 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR7_delayed) = 'X') and (TO_X01(WADDR7_previous) /= 'X')) then
             assert false
             report ": WADDR7 unknown"
             severity Warning;
            end if;
           else 
             RAM_di_int(7 downto 0) := DI7_delayed & DI6_delayed & DI5_delayed & DI4_delayed & DI3_delayed & DI2_delayed & DI1_delayed & DI0_delayed;
             memory_array(WADDR)  := RAM_di_int;
           end if;

         when others =>
          if (TO_X01(WBint_previous) /= 'X') then
             assert false
             report ": WRB or WBLKB unknown"
             severity Warning;
           end if;
      end case;
    end if;


 -----------------------------------------------------------
 --  Read Functional Section                              --
 -----------------------------------------------------------


    if (TO_X01(RCLKS_ipd) = 'X') then
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          RPE_zd := 'X';
       if (TO_X01(RCLKS_previous) /= 'X') then
         assert false
         report ": RCLK unknown"
         severity Warning;
       end if;
    elsif(RCLKS_ipd'event and RCLKS_ipd = '1') then

      case TO_X01(RBint_delayed) is
          when '1' =>
           null;
          when '0' =>

          if(RADDR < 0) then 
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          RPE_zd := 'X';
          if(TO_X01(RADDR0_delayed) = 'X') and (TO_X01(RADDR0_previous) /= 'X') then
             assert false
             report ": RADDR0 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR1_delayed) = 'X') and (TO_X01(RADDR1_previous) /= 'X') then
             assert false
             report ": RADDR1 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR2_delayed) = 'X') and (TO_X01(RADDR2_previous) /= 'X') then
             assert false
             report ": RADDR2 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR3_delayed) = 'X') and (TO_X01(RADDR3_previous) /= 'X') then
             assert false
             report ": RADDR3 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR4_delayed) = 'X') and (TO_X01(RADDR4_previous) /= 'X') then
             assert false
             report ": RADDR4 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR5_delayed) = 'X') and (TO_X01(RADDR5_previous) /= 'X') then
             assert false
             report ": RADDR5 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR6_delayed) = 'X') and (TO_X01(RADDR6_previous) /= 'X') then
             assert false
             report ": RADDR6 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR7_delayed) = 'X') and (TO_X01(RADDR7_previous) /= 'X') then
             assert false
             report ": RADDR7 unknown"
             severity Warning;
          end if;
          else  
            DO0_zd := memory_array(RADDR)(0);
            DO1_zd := memory_array(RADDR)(1);
            DO2_zd := memory_array(RADDR)(2);
            DO3_zd := memory_array(RADDR)(3);
            DO4_zd := memory_array(RADDR)(4);
            DO5_zd := memory_array(RADDR)(5);
            DO6_zd := memory_array(RADDR)(6);
            DO7_zd := memory_array(RADDR)(7);
            DO8_zd := memory_array(RADDR)(8);
            do_par  := DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR DO3_zd XOR DO2_zd XOR DO1_zd XOR DO0_zd;
            par_f <= do_par;
            if (do_par = 'X') then
              RPE_zd := 'X';
            elsif ( TO_X01 ( PARODD_delayed ) = 'X' ) then
              RPE_zd := 'X';
            else
              if ( do_par /= PARODD_delayed ) then
                RPE_zd  :=  '1';
              else
                RPE_zd  :=  '0';
              end if;
            end if;
        end if;

         when others =>
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          RPE_zd := 'X';
          if(TO_X01(RBint_previous) /= 'X') then
             assert false
             report ": RDB or RBLKB unknown "
             severity Warning;
           end if;
         end case;
       end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       WCLKS_previous  := WCLKS_ipd;
       RCLKS_previous  := RCLKS_ipd;
       RBint_previous := RBint_delayed;
       RBint_delayed  := RBint;
       WBint_previous  := WBint_delayed;
       WBint_delayed   := WBint;
       DI0_delayed     := DI0_ipd;
       DI1_delayed     := DI1_ipd;
       DI2_delayed     := DI2_ipd;
       DI3_delayed     := DI3_ipd;
       DI4_delayed     := DI4_ipd;
       DI5_delayed     := DI5_ipd;
       DI6_delayed     := DI6_ipd;
       DI7_delayed     := DI7_ipd;
       DI8_delayed     := DI8_ipd;
       RADDR0_previous := RADDR0_delayed;
       RADDR0_delayed  := RADDR0_ipd;
       RADDR1_previous := RADDR1_delayed;
       RADDR1_delayed  := RADDR1_ipd;
       RADDR2_previous := RADDR2_delayed;
       RADDR2_delayed  := RADDR2_ipd;
       RADDR3_previous := RADDR3_delayed;
       RADDR3_delayed  := RADDR3_ipd;
       RADDR4_previous := RADDR4_delayed;
       RADDR4_delayed  := RADDR4_ipd;
       RADDR5_previous := RADDR5_delayed;
       RADDR5_delayed  := RADDR5_ipd;
       RADDR6_previous := RADDR6_delayed;
       RADDR6_delayed  := RADDR6_ipd;
       RADDR7_previous := RADDR7_delayed;
       RADDR7_delayed  := RADDR7_ipd;
       WADDR0_previous := WADDR0_delayed;
       WADDR0_delayed  := WADDR0_ipd;
       WADDR1_previous := WADDR1_delayed;
       WADDR1_delayed  := WADDR1_ipd;
       WADDR2_previous := WADDR2_delayed;
       WADDR2_delayed  := WADDR2_ipd;
       WADDR3_previous := WADDR3_delayed;
       WADDR3_delayed  := WADDR3_ipd;
       WADDR4_previous := WADDR4_delayed;
       WADDR4_delayed  := WADDR4_ipd;
       WADDR5_previous := WADDR5_delayed;
       WADDR5_delayed  := WADDR5_ipd;
       WADDR6_previous := WADDR6_delayed;
       WADDR6_delayed  := WADDR6_ipd;
       WADDR7_previous := WADDR7_delayed;
       WADDR7_delayed  := WADDR7_ipd;
       PARODD_previous := PARODD_delayed; 
       PARODD_delayed  := PARODD_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
           OutSignal     => DOS,
           GlitchData    => DOS_GlitchData,
           OutSignalName => "DOS",
           OutTemp       => DOS_zd,
           Paths  =>  (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),
           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
             OutSignal     => WPE,
             GlitchData    => WPE_GlitchData,
             OutSignalName => "WPE",
             OutTemp       => WPE_zd,
             Paths =>   (0 => (WCLKS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_WCLKS_WPE), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
         OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => RPE,
           GlitchData    => RPE_GlitchData,
           OutSignalName => "RPE",
           OutTemp       => RPE_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_RPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
LIBRARY STD;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

USE std.textio.all;
USE ieee.std_logic_textio.all;
LIBRARY a500k;
USE a500k.all;

entity RAM256x9SSTP is 

   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tpw_WCLKS_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                           : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 7.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   WCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');

ATTRIBUTE VITAL_LEVEL0 OF RAM256x9SSTP : entity IS True ;
END RAM256x9SSTP;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of RAM256x9SSTP is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal WADDR0_ipd : std_ulogic := 'X';
   signal WADDR1_ipd : std_ulogic := 'X';
   signal WADDR2_ipd : std_ulogic := 'X';
   signal WADDR3_ipd : std_ulogic := 'X';
   signal WADDR4_ipd : std_ulogic := 'X';
   signal WADDR5_ipd : std_ulogic := 'X';
   signal WADDR6_ipd : std_ulogic := 'X';
   signal WADDR7_ipd : std_ulogic := 'X';
   signal RADDR0_ipd : std_ulogic := 'X';
   signal RADDR1_ipd : std_ulogic := 'X';
   signal RADDR2_ipd : std_ulogic := 'X';
   signal RADDR3_ipd : std_ulogic := 'X';
   signal RADDR4_ipd : std_ulogic := 'X';
   signal RADDR5_ipd : std_ulogic := 'X';
   signal RADDR6_ipd : std_ulogic := 'X';
   signal RADDR7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal WCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

	-- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';
   signal INIT_MEM   : std_logic:= '0';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic:= 'X';
   signal par_f2     : std_logic:= 'X';

 begin  --  VITAL_ACT
   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (WADDR0_ipd, WADDR0, VitalExtendToFillDelay(tipd_WADDR0));
   VitalWireDelay (WADDR1_ipd, WADDR1, VitalExtendToFillDelay(tipd_WADDR1));
   VitalWireDelay (WADDR2_ipd, WADDR2, VitalExtendToFillDelay(tipd_WADDR2));
   VitalWireDelay (WADDR3_ipd, WADDR3, VitalExtendToFillDelay(tipd_WADDR3));
   VitalWireDelay (WADDR4_ipd, WADDR4, VitalExtendToFillDelay(tipd_WADDR4));
   VitalWireDelay (WADDR5_ipd, WADDR5, VitalExtendToFillDelay(tipd_WADDR5));
   VitalWireDelay (WADDR6_ipd, WADDR6, VitalExtendToFillDelay(tipd_WADDR6));
   VitalWireDelay (WADDR7_ipd, WADDR7, VitalExtendToFillDelay(tipd_WADDR7));
   VitalWireDelay (RADDR0_ipd, RADDR0, VitalExtendToFillDelay(tipd_RADDR0));
   VitalWireDelay (RADDR1_ipd, RADDR1, VitalExtendToFillDelay(tipd_RADDR1));
   VitalWireDelay (RADDR2_ipd, RADDR2, VitalExtendToFillDelay(tipd_RADDR2));
   VitalWireDelay (RADDR3_ipd, RADDR3, VitalExtendToFillDelay(tipd_RADDR3));
   VitalWireDelay (RADDR4_ipd, RADDR4, VitalExtendToFillDelay(tipd_RADDR4));
   VitalWireDelay (RADDR5_ipd, RADDR5, VitalExtendToFillDelay(tipd_RADDR5));
   VitalWireDelay (RADDR6_ipd, RADDR6, VitalExtendToFillDelay(tipd_RADDR6));
   VitalWireDelay (RADDR7_ipd, RADDR7, VitalExtendToFillDelay(tipd_RADDR7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (WCLKS_ipd, WCLKS, VitalExtendToFillDelay(tipd_WCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

---------------------------------------------------------------
--                  Behavior Section                         --
---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);


    PROCESS
    BEGIN
      INIT_MEM <= '1';
      WAIT;
    END PROCESS;

    VITALBehavior : process (INIT_MEM, 
                          RADDR0_ipd, RADDR1_ipd, RADDR2_ipd, RADDR3_ipd, RADDR4_ipd, RADDR5_ipd, RADDR6_ipd, RADDR7_ipd, 
                          WADDR0_ipd, WADDR1_ipd, WADDR2_ipd, WADDR3_ipd, WADDR4_ipd, WADDR5_ipd, WADDR6_ipd, WADDR7_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd 
                          )

    -- some internal veriable declaration
     variable RAM_di_int         : std_logic_vector(8 downto 0);
     variable memory_array       : MEM_TYPE := (others =>(others => 'X'));
     variable do_par             : std_logic:= 'X';
     variable tmp_par            : std_logic:= 'X';
     variable tmp_par2           : std_logic:= 'X';
     variable wpe_var            : std_logic:= 'X';

     --  Read Timing Check Results
     variable Tviol_RADDR0_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR0_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR1_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR2_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR3_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR4_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR5_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR6_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR7_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable Tviol_WADDR0_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR0_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR1_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR2_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR3_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR4_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR5_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR6_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR7_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI0_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI1_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI2_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI3_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI4_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI5_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI6_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI7_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI8_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_WCLKS_posedge    : X01                 := '0';
     variable TmDt_WRB_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_WCLKS_posedge  : X01                 := '0';
     variable TmDt_WBLKB_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WCLKS                : X01                 := '0';
     variable Tviol_WCLKS_RCLKS_posedge  : X01                 := '0';
     variable TmDt_WCLKS_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results

     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     variable DO0_zd : std_ulogic;
     variable DO1_zd : std_ulogic;
     variable DO2_zd : std_ulogic;
     variable DO3_zd : std_ulogic;
     variable DO4_zd : std_ulogic;
     variable DO5_zd : std_ulogic;
     variable DO6_zd : std_ulogic;
     variable DO7_zd : std_ulogic;
     variable DO8_zd : std_ulogic;
     variable RPE_zd : std_ulogic;
     variable WPE_zd : std_ulogic;
     variable DOS_zd : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData  : VitalGlitchDataType;
     variable DO1_GlitchData  : VitalGlitchDataType;
     variable DO2_GlitchData  : VitalGlitchDataType;
     variable DO3_GlitchData  : VitalGlitchDataType;
     variable DO4_GlitchData  : VitalGlitchDataType;
     variable DO5_GlitchData  : VitalGlitchDataType;
     variable DO6_GlitchData  : VitalGlitchDataType;
     variable DO7_GlitchData  : VitalGlitchDataType;
     variable DO8_GlitchData  : VitalGlitchDataType;
     variable DOS_GlitchData  : VitalGlitchDataType;

     -- last value variables
     variable WCLKS_previous  : std_ulogic := 'X';
     variable RCLKS_previous  : std_ulogic := 'X';
     variable RBint_delayed   : std_ulogic := 'X';
     variable RBint_previous  : std_ulogic := 'X';
     variable WBint_delayed   : std_ulogic := 'X';
     variable WBint_previous  : std_ulogic := 'X';
     variable DIS_previous    : std_ulogic := 'X';
     variable DI0_delayed     : std_ulogic := 'X';
     variable DI1_delayed     : std_ulogic := 'X';
     variable DI2_delayed     : std_ulogic := 'X';
     variable DI3_delayed     : std_ulogic := 'X';
     variable DI4_delayed     : std_ulogic := 'X';
     variable DI5_delayed     : std_ulogic := 'X';
     variable DI6_delayed     : std_ulogic := 'X';
     variable DI7_delayed     : std_ulogic := 'X';
     variable DI8_delayed     : std_ulogic := 'X';
     variable RADDR0_delayed  : std_ulogic := 'X';
     variable RADDR1_delayed  : std_ulogic := 'X';
     variable RADDR2_delayed  : std_ulogic := 'X';
     variable RADDR3_delayed  : std_ulogic := 'X';
     variable RADDR4_delayed  : std_ulogic := 'X';
     variable RADDR5_delayed  : std_ulogic := 'X';
     variable RADDR6_delayed  : std_ulogic := 'X';
     variable RADDR7_delayed  : std_ulogic := 'X';
     variable RADDR0_previous : std_ulogic := 'X';
     variable RADDR1_previous : std_ulogic := 'X';
     variable RADDR2_previous : std_ulogic := 'X';
     variable RADDR3_previous : std_ulogic := 'X';
     variable RADDR4_previous : std_ulogic := 'X';
     variable RADDR5_previous : std_ulogic := 'X';
     variable RADDR6_previous : std_ulogic := 'X';
     variable RADDR7_previous : std_ulogic := 'X';
     variable WADDR0_delayed  : std_ulogic := 'X';
     variable WADDR1_delayed  : std_ulogic := 'X';
     variable WADDR2_delayed  : std_ulogic := 'X';
     variable WADDR3_delayed  : std_ulogic := 'X';
     variable WADDR4_delayed  : std_ulogic := 'X';
     variable WADDR5_delayed  : std_ulogic := 'X';
     variable WADDR6_delayed  : std_ulogic := 'X';
     variable WADDR7_delayed  : std_ulogic := 'X';
     variable WADDR0_previous : std_ulogic := 'X';
     variable WADDR1_previous : std_ulogic := 'X';
     variable WADDR2_previous : std_ulogic := 'X';
     variable WADDR3_previous : std_ulogic := 'X';
     variable WADDR4_previous : std_ulogic := 'X';
     variable WADDR5_previous : std_ulogic := 'X';
     variable WADDR6_previous : std_ulogic := 'X';
     variable WADDR7_previous : std_ulogic := 'X';

     variable PARODD_delayed  : std_ulogic := 'X';
     variable PARODD_previous : std_ulogic := 'X';

     variable inline    : LINE;
     variable indata    : std_logic_vector(8 downto 0);
     variable resdata   : std_logic_vector(8 downto 0);
     variable i         : integer:=0;
     file     memfile   : text;
     variable status         : file_open_status;

 begin -- process VITALBehavior

  -----------------------------------------------------------
  --    Initialize memory file from MEMORYFILE string      --
  -----------------------------------------------------------


  if ( INIT_MEM'EVENT and INIT_MEM = '1') then
    file_open(status, memfile, MEMORYFILE, read_mode);
    if ( status=open_ok ) then
      while((i < 256) and (not ENDFILE(memfile))) loop
        readline(memfile,inline);
        read(inline,indata);
        resdata := indata;
        memory_array(i) := resdata;
        i := i+1;
      end loop;
    else
      assert ( MEMORYFILE'length = 0 )
        report "Failed to open RAM256x9SSTP memory initialization file in read mode"
        severity Note;
    end if;
    file_close(memfile);
  end if;


     if (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      WADDR := ((INT(WADDR7_delayed)*128)+(INT(WADDR6_delayed)*64)+(INT(
               WADDR5_delayed)*32) + (INT(WADDR4_delayed)*16) + 
               (INT(WADDR3_delayed)*8) + (INT(WADDR2_delayed)*4) + (INT(
               WADDR1_delayed)*2) + (INT(WADDR0_delayed)*1));
     end if;

   -- Convert Read Address Signal to Integer
     if (RCLKS_ipd'EVENT AND RCLKS_ipd = '1') then
      RADDR := ((INT(RADDR7_delayed)*128)+(INT(RADDR6_delayed)*64)+(INT(
               RADDR5_delayed)*32) + (INT(RADDR4_delayed)*16) + 
               (INT(RADDR3_delayed)*8) + (INT(RADDR2_delayed)*4) + (INT(
               RADDR1_delayed)*2) + (INT(RADDR0_delayed)*1));
     end if;

if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

 -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SSTP",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_WADDR0_WCLKS_posedge,
                             TmDt_WADDR0_WCLKS_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR0_WCLKS_posedge_posedge,
                             tsetup_WADDR0_WCLKS_posedge_posedge,
                             thold_WADDR0_WCLKS_posedge_posedge,
                             thold_WADDR0_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WCLKS_posedge,
                             TmDt_WADDR0_WCLKS_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR0_WCLKS_negedge_posedge,
                             tsetup_WADDR0_WCLKS_negedge_posedge,
                             thold_WADDR0_WCLKS_negedge_posedge,
                             thold_WADDR0_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WCLKS_posedge,
                             TmDt_WADDR1_WCLKS_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR1_WCLKS_posedge_posedge,
                             tsetup_WADDR1_WCLKS_posedge_posedge,
                             thold_WADDR1_WCLKS_posedge_posedge,
                             thold_WADDR1_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WCLKS_posedge,
                             TmDt_WADDR1_WCLKS_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR1_WCLKS_negedge_posedge,
                             tsetup_WADDR1_WCLKS_negedge_posedge,
                             thold_WADDR1_WCLKS_negedge_posedge,
                             thold_WADDR1_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WCLKS_posedge,
                             TmDt_WADDR2_WCLKS_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR2_WCLKS_posedge_posedge,
                             tsetup_WADDR2_WCLKS_posedge_posedge,
                             thold_WADDR2_WCLKS_posedge_posedge,
                             thold_WADDR2_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WCLKS_posedge,
                             TmDt_WADDR2_WCLKS_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR2_WCLKS_negedge_posedge,
                             tsetup_WADDR2_WCLKS_negedge_posedge,
                             thold_WADDR2_WCLKS_negedge_posedge,
                             thold_WADDR2_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WCLKS_posedge,
                             TmDt_WADDR3_WCLKS_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR3_WCLKS_posedge_posedge,
                             tsetup_WADDR3_WCLKS_posedge_posedge,
                             thold_WADDR3_WCLKS_posedge_posedge,
                             thold_WADDR3_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WCLKS_posedge,
                             TmDt_WADDR3_WCLKS_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR3_WCLKS_negedge_posedge,
                             tsetup_WADDR3_WCLKS_negedge_posedge,
                             thold_WADDR3_WCLKS_negedge_posedge,
                             thold_WADDR3_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WCLKS_posedge,
                             TmDt_WADDR4_WCLKS_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR4_WCLKS_posedge_posedge,
                             tsetup_WADDR4_WCLKS_posedge_posedge,
                             thold_WADDR4_WCLKS_posedge_posedge,
                             thold_WADDR4_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WCLKS_posedge,
                             TmDt_WADDR4_WCLKS_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR4_WCLKS_negedge_posedge,
                             tsetup_WADDR4_WCLKS_negedge_posedge,
                             thold_WADDR4_WCLKS_negedge_posedge,
                             thold_WADDR4_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WCLKS_posedge,
                             TmDt_WADDR5_WCLKS_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR5_WCLKS_posedge_posedge,
                             tsetup_WADDR5_WCLKS_posedge_posedge,
                             thold_WADDR5_WCLKS_posedge_posedge,
                             thold_WADDR5_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WCLKS_posedge,
                             TmDt_WADDR5_WCLKS_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR5_WCLKS_negedge_posedge,
                             tsetup_WADDR5_WCLKS_negedge_posedge,
                             thold_WADDR5_WCLKS_negedge_posedge,
                             thold_WADDR5_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WCLKS_posedge,
                             TmDt_WADDR6_WCLKS_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR6_WCLKS_posedge_posedge,
                             tsetup_WADDR6_WCLKS_posedge_posedge,
                             thold_WADDR6_WCLKS_posedge_posedge,
                             thold_WADDR6_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WCLKS_posedge,
                             TmDt_WADDR6_WCLKS_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR6_WCLKS_negedge_posedge,
                             tsetup_WADDR6_WCLKS_negedge_posedge,
                             thold_WADDR6_WCLKS_negedge_posedge,
                             thold_WADDR6_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WCLKS_posedge,
                             TmDt_WADDR7_WCLKS_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR7_WCLKS_posedge_posedge,
                             tsetup_WADDR7_WCLKS_posedge_posedge,
                             thold_WADDR7_WCLKS_posedge_posedge,
                             thold_WADDR7_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WCLKS_posedge,
                             TmDt_WADDR7_WCLKS_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR7_WCLKS_negedge_posedge,
                             tsetup_WADDR7_WCLKS_negedge_posedge,
                             thold_WADDR7_WCLKS_negedge_posedge,
                             thold_WADDR7_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_posedge_posedge,
                             tsetup_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_negedge_posedge,
                             tsetup_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_posedge_posedge,
                             tsetup_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_negedge_posedge,
                             tsetup_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_posedge_posedge,
                             tsetup_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_negedge_posedge,
                             tsetup_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_posedge_posedge,
                             tsetup_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_negedge_posedge,
                             tsetup_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_posedge_posedge,
                             tsetup_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_negedge_posedge,
                             tsetup_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_posedge_posedge,
                             tsetup_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_negedge_posedge,
                             tsetup_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_posedge_posedge,
                             tsetup_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_negedge_posedge,
                             tsetup_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_posedge_posedge,
                             tsetup_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_negedge_posedge,
                             tsetup_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_posedge_posedge,
                             tsetup_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_negedge_posedge,
                             tsetup_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

 -- setup hold WEN, WBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_posedge_posedge,
                             tsetup_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_negedge_posedge,
                             tsetup_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

  --   Period of WCLK
      VitalPeriodPulseCheck ( Pviol_WCLKS,
                              PeriodData_WCLKS,
                              WCLKS_ipd, "WCLKS",
                              0.0 ns,
                              tperiod_WCLKS,
                              tpw_WCLKS_posedge,
                              tpw_WCLKS_negedge,
                              (To_X01(WBLKB_ipd) = '0') AND (To_X01(WRB_ipd) = '0'),
                             InstancePath & "/RAM256x9SSTP",
                              True,
                              True,
                              WARNING
                              );
   ------------------------------------------------------------
   --        Timing Checking for Read and write conflict     --
   ------------------------------------------------------------
       VitalSetupHoldCheck ( Tviol_WCLKS_RCLKS_posedge,
                             TmDt_WCLKS_RCLKS_posedge,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_WCLKS_RCLKS_posedge_posedge,
                             0.0 ns,
                             thold_WCLKS_RCLKS_posedge_posedge,
                             0.0 ns,
                             (To_X01(RBint) = '0') AND (To_X01(WBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

 end if;

   ------------------------------------------------------------
   --         WPE generating  block                            -
   ------------------------------------------------------------

     if (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
        tmp_par  := DI7_delayed XOR DI6_delayed XOR DI5_delayed XOR DI4_delayed XOR DI3_delayed XOR DI2_delayed XOR DI1_delayed XOR DI0_delayed;
        if (tmp_par   /= PARODD_delayed) then
           wpe_var     :=  '1';
        else
           wpe_var     :=  '0';
        end if;
        RAM_di_int(8) := wpe_var;
        WPE_zd := wpe_var;
     end if;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

    if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
    end if; 

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

  if (TO_X01(WCLKS_ipd)='X') then
   if (TO_X01(WCLKS_previous) /= 'X') then
    assert false
    report ": WCLK unknown"
    severity Warning;
    end if;
   elsif (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      case TO_X01(WBint_delayed) is
          when '1' =>
            null;
          when '0' =>
           if(WADDR < 0) then
            if ((TO_X01(WADDR0_delayed) = 'X') and (TO_X01(WADDR0_previous) /= 'X')) then
             assert false
             report ": WADDR0 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR1_delayed) = 'X') and (TO_X01(WADDR1_previous) /= 'X')) then
             assert false
             report ": WADDR1 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR2_delayed) = 'X') and (TO_X01(WADDR2_previous) /= 'X')) then
             assert false
             report ": WADDR2 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR3_delayed) = 'X') and (TO_X01(WADDR3_previous) /= 'X')) then
             assert false
             report ": WADDR3 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR4_delayed) = 'X') and (TO_X01(WADDR4_previous) /= 'X')) then
             assert false
             report ": WADDR4 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR5_delayed) = 'X') and (TO_X01(WADDR5_previous) /= 'X')) then
             assert false
             report ": WADDR5 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR6_delayed) = 'X') and (TO_X01(WADDR6_previous) /= 'X')) then
             assert false
             report ": WADDR6 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR7_delayed) = 'X') and (TO_X01(WADDR7_previous) /= 'X')) then
             assert false
             report ": WADDR7 unknown"
             severity Warning;
            end if;
           else 
             RAM_di_int(7 downto 0) := DI7_delayed & DI6_delayed & DI5_delayed & DI4_delayed & DI3_delayed & DI2_delayed & DI1_delayed & DI0_delayed;
             memory_array(WADDR)  := RAM_di_int;
           end if;

         when others =>
          if (TO_X01(WBint_previous) /= 'X') then
             assert false
             report ": WRB or WBLKB unknown"
             severity Warning;
           end if;
      end case;
    end if;


 -----------------------------------------------------------
 --  Read Functional Section                              --
 -----------------------------------------------------------


    if (TO_X01(RCLKS_ipd) = 'X') then
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          RPE_zd := 'X';
       if (TO_X01(RCLKS_previous) /= 'X') then
         assert false
         report ": RCLK unknown"
         severity Warning;
       end if;
    elsif(RCLKS_ipd'event and RCLKS_ipd = '1') then

      case TO_X01(RBint_delayed) is
          when '1' =>
           null;
          when '0' =>

          if(RADDR < 0) then 
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          if(TO_X01(RADDR0_delayed) = 'X') and (TO_X01(RADDR0_previous) /= 'X') then
             assert false
             report ": RADDR0 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR1_delayed) = 'X') and (TO_X01(RADDR1_previous) /= 'X') then
             assert false
             report ": RADDR1 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR2_delayed) = 'X') and (TO_X01(RADDR2_previous) /= 'X') then
             assert false
             report ": RADDR2 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR3_delayed) = 'X') and (TO_X01(RADDR3_previous) /= 'X') then
             assert false
             report ": RADDR3 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR4_delayed) = 'X') and (TO_X01(RADDR4_previous) /= 'X') then
             assert false
             report ": RADDR4 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR5_delayed) = 'X') and (TO_X01(RADDR5_previous) /= 'X') then
             assert false
             report ": RADDR5 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR6_delayed) = 'X') and (TO_X01(RADDR6_previous) /= 'X') then
             assert false
             report ": RADDR6 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR7_delayed) = 'X') and (TO_X01(RADDR7_previous) /= 'X') then
             assert false
             report ": RADDR7 unknown"
             severity Warning;
          end if;
          else  
            DO0_zd := memory_array(RADDR)(0);
            DO1_zd := memory_array(RADDR)(1);
            DO2_zd := memory_array(RADDR)(2);
            DO3_zd := memory_array(RADDR)(3);
            DO4_zd := memory_array(RADDR)(4);
            DO5_zd := memory_array(RADDR)(5);
            DO6_zd := memory_array(RADDR)(6);
            DO7_zd := memory_array(RADDR)(7);
            DO8_zd := memory_array(RADDR)(8);
        end if;

         when others =>
          DO0_zd := 'X';
          DO1_zd := 'X';
          DO2_zd := 'X';
          DO3_zd := 'X';
          DO4_zd := 'X';
          DO5_zd := 'X';
          DO6_zd := 'X';
          DO7_zd := 'X';
          DO8_zd := 'X';
          if(TO_X01(RBint_previous) /= 'X') then
             assert false
             report ": RDB or RBLKB unknown "
             severity Warning;
           end if;
         end case;
       end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       WCLKS_previous  := WCLKS_ipd;
       RCLKS_previous  := RCLKS_ipd;
       RBint_previous := RBint_delayed;
       RBint_delayed  := RBint;
       WBint_previous  := WBint_delayed;
       WBint_delayed   := WBint;
       DI0_delayed     := DI0_ipd;
       DI1_delayed     := DI1_ipd;
       DI2_delayed     := DI2_ipd;
       DI3_delayed     := DI3_ipd;
       DI4_delayed     := DI4_ipd;
       DI5_delayed     := DI5_ipd;
       DI6_delayed     := DI6_ipd;
       DI7_delayed     := DI7_ipd;
       DI8_delayed     := DI8_ipd;
       RADDR0_previous := RADDR0_delayed;
       RADDR0_delayed  := RADDR0_ipd;
       RADDR1_previous := RADDR1_delayed;
       RADDR1_delayed  := RADDR1_ipd;
       RADDR2_previous := RADDR2_delayed;
       RADDR2_delayed  := RADDR2_ipd;
       RADDR3_previous := RADDR3_delayed;
       RADDR3_delayed  := RADDR3_ipd;
       RADDR4_previous := RADDR4_delayed;
       RADDR4_delayed  := RADDR4_ipd;
       RADDR5_previous := RADDR5_delayed;
       RADDR5_delayed  := RADDR5_ipd;
       RADDR6_previous := RADDR6_delayed;
       RADDR6_delayed  := RADDR6_ipd;
       RADDR7_previous := RADDR7_delayed;
       RADDR7_delayed  := RADDR7_ipd;
       WADDR0_previous := WADDR0_delayed;
       WADDR0_delayed  := WADDR0_ipd;
       WADDR1_previous := WADDR1_delayed;
       WADDR1_delayed  := WADDR1_ipd;
       WADDR2_previous := WADDR2_delayed;
       WADDR2_delayed  := WADDR2_ipd;
       WADDR3_previous := WADDR3_delayed;
       WADDR3_delayed  := WADDR3_ipd;
       WADDR4_previous := WADDR4_delayed;
       WADDR4_delayed  := WADDR4_ipd;
       WADDR5_previous := WADDR5_delayed;
       WADDR5_delayed  := WADDR5_ipd;
       WADDR6_previous := WADDR6_delayed;
       WADDR6_delayed  := WADDR6_ipd;
       WADDR7_previous := WADDR7_delayed;
       WADDR7_delayed  := WADDR7_ipd;
       PARODD_previous := PARODD_delayed; 
       PARODD_delayed  := PARODD_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
           OutSignal     => DOS,
           GlitchData    => DOS_GlitchData,
           OutSignalName => "DOS",
           OutTemp       => DOS_zd,
           Paths  =>  (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),
           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
LIBRARY STD;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

USE std.textio.all;
USE ieee.std_logic_textio.all;
LIBRARY a500k;
USE a500k.all;

entity RAM256x9SSR is 

   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_WCLKS_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tpw_WCLKS_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                           : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 7.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';
   WPE    :  OUT STD_LOGIC := 'X';
   RPE    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   WCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');

ATTRIBUTE VITAL_LEVEL0 OF RAM256x9SSR : entity IS True ;
END RAM256x9SSR;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of RAM256x9SSR is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal WADDR0_ipd : std_ulogic := 'X';
   signal WADDR1_ipd : std_ulogic := 'X';
   signal WADDR2_ipd : std_ulogic := 'X';
   signal WADDR3_ipd : std_ulogic := 'X';
   signal WADDR4_ipd : std_ulogic := 'X';
   signal WADDR5_ipd : std_ulogic := 'X';
   signal WADDR6_ipd : std_ulogic := 'X';
   signal WADDR7_ipd : std_ulogic := 'X';
   signal RADDR0_ipd : std_ulogic := 'X';
   signal RADDR1_ipd : std_ulogic := 'X';
   signal RADDR2_ipd : std_ulogic := 'X';
   signal RADDR3_ipd : std_ulogic := 'X';
   signal RADDR4_ipd : std_ulogic := 'X';
   signal RADDR5_ipd : std_ulogic := 'X';
   signal RADDR6_ipd : std_ulogic := 'X';
   signal RADDR7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal WCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

	-- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';
   signal INIT_MEM   : std_logic:= '0';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic:= 'X';
   signal par_f2     : std_logic:= 'X';

 begin  --  VITAL_ACT
   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (WADDR0_ipd, WADDR0, VitalExtendToFillDelay(tipd_WADDR0));
   VitalWireDelay (WADDR1_ipd, WADDR1, VitalExtendToFillDelay(tipd_WADDR1));
   VitalWireDelay (WADDR2_ipd, WADDR2, VitalExtendToFillDelay(tipd_WADDR2));
   VitalWireDelay (WADDR3_ipd, WADDR3, VitalExtendToFillDelay(tipd_WADDR3));
   VitalWireDelay (WADDR4_ipd, WADDR4, VitalExtendToFillDelay(tipd_WADDR4));
   VitalWireDelay (WADDR5_ipd, WADDR5, VitalExtendToFillDelay(tipd_WADDR5));
   VitalWireDelay (WADDR6_ipd, WADDR6, VitalExtendToFillDelay(tipd_WADDR6));
   VitalWireDelay (WADDR7_ipd, WADDR7, VitalExtendToFillDelay(tipd_WADDR7));
   VitalWireDelay (RADDR0_ipd, RADDR0, VitalExtendToFillDelay(tipd_RADDR0));
   VitalWireDelay (RADDR1_ipd, RADDR1, VitalExtendToFillDelay(tipd_RADDR1));
   VitalWireDelay (RADDR2_ipd, RADDR2, VitalExtendToFillDelay(tipd_RADDR2));
   VitalWireDelay (RADDR3_ipd, RADDR3, VitalExtendToFillDelay(tipd_RADDR3));
   VitalWireDelay (RADDR4_ipd, RADDR4, VitalExtendToFillDelay(tipd_RADDR4));
   VitalWireDelay (RADDR5_ipd, RADDR5, VitalExtendToFillDelay(tipd_RADDR5));
   VitalWireDelay (RADDR6_ipd, RADDR6, VitalExtendToFillDelay(tipd_RADDR6));
   VitalWireDelay (RADDR7_ipd, RADDR7, VitalExtendToFillDelay(tipd_RADDR7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (WCLKS_ipd, WCLKS, VitalExtendToFillDelay(tipd_WCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

---------------------------------------------------------------
--                  Behavior Section                         --
---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);


    PROCESS
    BEGIN
      INIT_MEM <= '1';
      WAIT;
    END PROCESS;

    VITALBehavior : process (INIT_MEM, 
                          RADDR0_ipd, RADDR1_ipd, RADDR2_ipd, RADDR3_ipd, RADDR4_ipd, RADDR5_ipd, RADDR6_ipd, RADDR7_ipd, 
                          WADDR0_ipd, WADDR1_ipd, WADDR2_ipd, WADDR3_ipd, WADDR4_ipd, WADDR5_ipd, WADDR6_ipd, WADDR7_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd 
                          )

    -- some internal veriable declaration
     variable RAM_di_int         : std_logic_vector(8 downto 0);
     variable memory_array       : MEM_TYPE := (others =>(others => 'X'));
     variable do_par             : std_logic:= 'X';
     variable tmp_par            : std_logic:= 'X';
     variable tmp_par2           : std_logic:= 'X';
     variable wpe_var            : std_logic:= 'X';

     --  Read Timing Check Results
     variable Tviol_RADDR0_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR0_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR1_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR2_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR3_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR4_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR5_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR6_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR7_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable Tviol_WADDR0_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR0_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR1_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR2_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR3_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR4_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR5_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR6_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR7_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI0_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI1_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI2_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI3_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI4_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI5_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI6_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI7_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI8_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_WCLKS_posedge    : X01                 := '0';
     variable TmDt_WRB_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_WCLKS_posedge  : X01                 := '0';
     variable TmDt_WBLKB_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WCLKS                : X01                 := '0';
     variable Tviol_WCLKS_RCLKS_posedge  : X01                 := '0';
     variable TmDt_WCLKS_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results

     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     variable DO0_zd : std_ulogic;
     variable DO1_zd : std_ulogic;
     variable DO2_zd : std_ulogic;
     variable DO3_zd : std_ulogic;
     variable DO4_zd : std_ulogic;
     variable DO5_zd : std_ulogic;
     variable DO6_zd : std_ulogic;
     variable DO7_zd : std_ulogic;
     variable DO8_zd : std_ulogic;
     variable RPE_zd : std_ulogic;
     variable WPE_zd : std_ulogic;
     variable DOS_zd : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData  : VitalGlitchDataType;
     variable DO1_GlitchData  : VitalGlitchDataType;
     variable DO2_GlitchData  : VitalGlitchDataType;
     variable DO3_GlitchData  : VitalGlitchDataType;
     variable DO4_GlitchData  : VitalGlitchDataType;
     variable DO5_GlitchData  : VitalGlitchDataType;
     variable DO6_GlitchData  : VitalGlitchDataType;
     variable DO7_GlitchData  : VitalGlitchDataType;
     variable DO8_GlitchData  : VitalGlitchDataType;
     variable RPE_GlitchData  : VitalGlitchDataType;
     variable WPE_GlitchData  : VitalGlitchDataType;
     variable DOS_GlitchData  : VitalGlitchDataType;

     -- last value variables
     variable WCLKS_previous  : std_ulogic := 'X';
     variable RCLKS_previous  : std_ulogic := 'X';
     variable RBint_delayed   : std_ulogic := 'X';
     variable RBint_previous  : std_ulogic := 'X';
     variable WBint_delayed   : std_ulogic := 'X';
     variable WBint_previous  : std_ulogic := 'X';
     variable DIS_previous    : std_ulogic := 'X';
     variable DI0_delayed     : std_ulogic := 'X';
     variable DI1_delayed     : std_ulogic := 'X';
     variable DI2_delayed     : std_ulogic := 'X';
     variable DI3_delayed     : std_ulogic := 'X';
     variable DI4_delayed     : std_ulogic := 'X';
     variable DI5_delayed     : std_ulogic := 'X';
     variable DI6_delayed     : std_ulogic := 'X';
     variable DI7_delayed     : std_ulogic := 'X';
     variable DI8_delayed     : std_ulogic := 'X';
     variable RADDR0_delayed  : std_ulogic := 'X';
     variable RADDR1_delayed  : std_ulogic := 'X';
     variable RADDR2_delayed  : std_ulogic := 'X';
     variable RADDR3_delayed  : std_ulogic := 'X';
     variable RADDR4_delayed  : std_ulogic := 'X';
     variable RADDR5_delayed  : std_ulogic := 'X';
     variable RADDR6_delayed  : std_ulogic := 'X';
     variable RADDR7_delayed  : std_ulogic := 'X';
     variable RADDR0_previous : std_ulogic := 'X';
     variable RADDR1_previous : std_ulogic := 'X';
     variable RADDR2_previous : std_ulogic := 'X';
     variable RADDR3_previous : std_ulogic := 'X';
     variable RADDR4_previous : std_ulogic := 'X';
     variable RADDR5_previous : std_ulogic := 'X';
     variable RADDR6_previous : std_ulogic := 'X';
     variable RADDR7_previous : std_ulogic := 'X';
     variable WADDR0_delayed  : std_ulogic := 'X';
     variable WADDR1_delayed  : std_ulogic := 'X';
     variable WADDR2_delayed  : std_ulogic := 'X';
     variable WADDR3_delayed  : std_ulogic := 'X';
     variable WADDR4_delayed  : std_ulogic := 'X';
     variable WADDR5_delayed  : std_ulogic := 'X';
     variable WADDR6_delayed  : std_ulogic := 'X';
     variable WADDR7_delayed  : std_ulogic := 'X';
     variable WADDR0_previous : std_ulogic := 'X';
     variable WADDR1_previous : std_ulogic := 'X';
     variable WADDR2_previous : std_ulogic := 'X';
     variable WADDR3_previous : std_ulogic := 'X';
     variable WADDR4_previous : std_ulogic := 'X';
     variable WADDR5_previous : std_ulogic := 'X';
     variable WADDR6_previous : std_ulogic := 'X';
     variable WADDR7_previous : std_ulogic := 'X';

     --  Pipelined temporary results
    variable RPE_stg1        : std_ulogic := 'X';
    variable DO0_stg1        : std_ulogic := 'X';
    variable DO1_stg1        : std_ulogic := 'X';
    variable DO2_stg1        : std_ulogic := 'X';
    variable DO3_stg1        : std_ulogic := 'X';
    variable DO4_stg1        : std_ulogic := 'X';
    variable DO5_stg1        : std_ulogic := 'X';
    variable DO6_stg1        : std_ulogic := 'X';
    variable DO7_stg1        : std_ulogic := 'X';
    variable DO8_stg1        : std_ulogic := 'X';

    variable PARODD_delayed  : std_ulogic := 'X';
    variable PARODD_previous : std_ulogic := 'X';

    variable inline    : LINE;
    variable indata    : std_logic_vector(8 downto 0);
    variable resdata   : std_logic_vector(8 downto 0);
    variable i         : integer:=0;
    file     memfile   : text;
    variable status         : file_open_status;

 begin -- process VITALBehavior


  -----------------------------------------------------------
  --    Initialize memory file from MEMORYFILE string      --
  -----------------------------------------------------------


  if ( INIT_MEM'EVENT and INIT_MEM = '1') then
    file_open(status, memfile, MEMORYFILE, read_mode);
    if ( status=open_ok ) then
      while((i < 256) and (not ENDFILE(memfile))) loop
        readline(memfile,inline);
        read(inline,indata);
        resdata := indata;
        memory_array(i) := resdata;
        i := i+1;
      end loop;
    else
      assert ( MEMORYFILE'length = 0 )
        report "Failed to open RAM256x9SSR memory initialization file in read mode"
        severity Note;
    end if;
    file_close(memfile);
  end if;


     if (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      WADDR := ((INT(WADDR7_delayed)*128)+(INT(WADDR6_delayed)*64)+(INT(
               WADDR5_delayed)*32) + (INT(WADDR4_delayed)*16) + 
               (INT(WADDR3_delayed)*8) + (INT(WADDR2_delayed)*4) + (INT(
               WADDR1_delayed)*2) + (INT(WADDR0_delayed)*1));
     end if;

   -- Convert Read Address Signal to Integer
     if (RCLKS_ipd'EVENT AND RCLKS_ipd = '1') then
      RADDR := ((INT(RADDR7_delayed)*128)+(INT(RADDR6_delayed)*64)+(INT(
               RADDR5_delayed)*32) + (INT(RADDR4_delayed)*16) + 
               (INT(RADDR3_delayed)*8) + (INT(RADDR2_delayed)*4) + (INT(
               RADDR1_delayed)*2) + (INT(RADDR0_delayed)*1));
     end if;

if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

 -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SSR",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_WADDR0_WCLKS_posedge,
                             TmDt_WADDR0_WCLKS_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR0_WCLKS_posedge_posedge,
                             tsetup_WADDR0_WCLKS_posedge_posedge,
                             thold_WADDR0_WCLKS_posedge_posedge,
                             thold_WADDR0_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WCLKS_posedge,
                             TmDt_WADDR0_WCLKS_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR0_WCLKS_negedge_posedge,
                             tsetup_WADDR0_WCLKS_negedge_posedge,
                             thold_WADDR0_WCLKS_negedge_posedge,
                             thold_WADDR0_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WCLKS_posedge,
                             TmDt_WADDR1_WCLKS_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR1_WCLKS_posedge_posedge,
                             tsetup_WADDR1_WCLKS_posedge_posedge,
                             thold_WADDR1_WCLKS_posedge_posedge,
                             thold_WADDR1_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WCLKS_posedge,
                             TmDt_WADDR1_WCLKS_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR1_WCLKS_negedge_posedge,
                             tsetup_WADDR1_WCLKS_negedge_posedge,
                             thold_WADDR1_WCLKS_negedge_posedge,
                             thold_WADDR1_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WCLKS_posedge,
                             TmDt_WADDR2_WCLKS_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR2_WCLKS_posedge_posedge,
                             tsetup_WADDR2_WCLKS_posedge_posedge,
                             thold_WADDR2_WCLKS_posedge_posedge,
                             thold_WADDR2_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WCLKS_posedge,
                             TmDt_WADDR2_WCLKS_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR2_WCLKS_negedge_posedge,
                             tsetup_WADDR2_WCLKS_negedge_posedge,
                             thold_WADDR2_WCLKS_negedge_posedge,
                             thold_WADDR2_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WCLKS_posedge,
                             TmDt_WADDR3_WCLKS_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR3_WCLKS_posedge_posedge,
                             tsetup_WADDR3_WCLKS_posedge_posedge,
                             thold_WADDR3_WCLKS_posedge_posedge,
                             thold_WADDR3_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WCLKS_posedge,
                             TmDt_WADDR3_WCLKS_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR3_WCLKS_negedge_posedge,
                             tsetup_WADDR3_WCLKS_negedge_posedge,
                             thold_WADDR3_WCLKS_negedge_posedge,
                             thold_WADDR3_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WCLKS_posedge,
                             TmDt_WADDR4_WCLKS_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR4_WCLKS_posedge_posedge,
                             tsetup_WADDR4_WCLKS_posedge_posedge,
                             thold_WADDR4_WCLKS_posedge_posedge,
                             thold_WADDR4_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WCLKS_posedge,
                             TmDt_WADDR4_WCLKS_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR4_WCLKS_negedge_posedge,
                             tsetup_WADDR4_WCLKS_negedge_posedge,
                             thold_WADDR4_WCLKS_negedge_posedge,
                             thold_WADDR4_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WCLKS_posedge,
                             TmDt_WADDR5_WCLKS_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR5_WCLKS_posedge_posedge,
                             tsetup_WADDR5_WCLKS_posedge_posedge,
                             thold_WADDR5_WCLKS_posedge_posedge,
                             thold_WADDR5_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WCLKS_posedge,
                             TmDt_WADDR5_WCLKS_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR5_WCLKS_negedge_posedge,
                             tsetup_WADDR5_WCLKS_negedge_posedge,
                             thold_WADDR5_WCLKS_negedge_posedge,
                             thold_WADDR5_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WCLKS_posedge,
                             TmDt_WADDR6_WCLKS_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR6_WCLKS_posedge_posedge,
                             tsetup_WADDR6_WCLKS_posedge_posedge,
                             thold_WADDR6_WCLKS_posedge_posedge,
                             thold_WADDR6_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WCLKS_posedge,
                             TmDt_WADDR6_WCLKS_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR6_WCLKS_negedge_posedge,
                             tsetup_WADDR6_WCLKS_negedge_posedge,
                             thold_WADDR6_WCLKS_negedge_posedge,
                             thold_WADDR6_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WCLKS_posedge,
                             TmDt_WADDR7_WCLKS_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR7_WCLKS_posedge_posedge,
                             tsetup_WADDR7_WCLKS_posedge_posedge,
                             thold_WADDR7_WCLKS_posedge_posedge,
                             thold_WADDR7_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WCLKS_posedge,
                             TmDt_WADDR7_WCLKS_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR7_WCLKS_negedge_posedge,
                             tsetup_WADDR7_WCLKS_negedge_posedge,
                             thold_WADDR7_WCLKS_negedge_posedge,
                             thold_WADDR7_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_posedge_posedge,
                             tsetup_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_negedge_posedge,
                             tsetup_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_posedge_posedge,
                             tsetup_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_negedge_posedge,
                             tsetup_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_posedge_posedge,
                             tsetup_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_negedge_posedge,
                             tsetup_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_posedge_posedge,
                             tsetup_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_negedge_posedge,
                             tsetup_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_posedge_posedge,
                             tsetup_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_negedge_posedge,
                             tsetup_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_posedge_posedge,
                             tsetup_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_negedge_posedge,
                             tsetup_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_posedge_posedge,
                             tsetup_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_negedge_posedge,
                             tsetup_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_posedge_posedge,
                             tsetup_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_negedge_posedge,
                             tsetup_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_posedge_posedge,
                             tsetup_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_negedge_posedge,
                             tsetup_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

 -- setup hold WEN, WBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_posedge_posedge,
                             tsetup_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_negedge_posedge,
                             tsetup_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

  --   Period of WCLK
      VitalPeriodPulseCheck ( Pviol_WCLKS,
                              PeriodData_WCLKS,
                              WCLKS_ipd, "WCLKS",
                              0.0 ns,
                              tperiod_WCLKS,
                              tpw_WCLKS_posedge,
                              tpw_WCLKS_negedge,
                              (To_X01(WBLKB_ipd) = '0') AND (To_X01(WRB_ipd) = '0'),
                             InstancePath & "/RAM256x9SSR",
                              True,
                              True,
                              WARNING
                              );
   ------------------------------------------------------------
   --        Timing Checking for Read and write conflict     --
   ------------------------------------------------------------
       VitalSetupHoldCheck ( Tviol_WCLKS_RCLKS_posedge,
                             TmDt_WCLKS_RCLKS_posedge,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_WCLKS_RCLKS_posedge_posedge,
                             0.0 ns,
                             thold_WCLKS_RCLKS_posedge_posedge,
                             0.0 ns,
                             (To_X01(RBint) = '0') AND (To_X01(WBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SSR",
                             True,
                             True,
                             WARNING
                             );

 end if;

   ------------------------------------------------------------
   --    wpe output                                           -
   ------------------------------------------------------------

   if ( PARODD_ipd'EVENT ) then
     RPE_zd := not RPE_zd;
     RPE_stg1 := not RPE_stg1;
     WPE_zd := not WPE_zd;
   end if;

   ------------------------------------------------------------
   --         WPE checking  block                            -
   ------------------------------------------------------------

     if ( WCLKS_ipd'EVENT ) then
        tmp_par  := DI7_delayed XOR DI6_delayed XOR DI5_delayed XOR DI4_delayed XOR DI3_delayed XOR DI2_delayed XOR DI1_delayed XOR DI0_delayed;
        tmp_par2 := (tmp_par xor DI8_delayed);

      if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
          ( TO_X01 ( WCLKS_ipd  ) = 'X' ) or 
          ( TO_X01 ( DI8_ipd )    = 'X' ) or
          ( TO_X01 ( DI7_ipd )    = 'X' ) or
          ( TO_X01 ( DI6_ipd )    = 'X' ) or
          ( TO_X01 ( DI5_ipd )    = 'X' ) or
          ( TO_X01 ( DI4_ipd )    = 'X' ) or
          ( TO_X01 ( DI3_ipd )    = 'X' ) or
          ( TO_X01 ( DI2_ipd )    = 'X' ) or
          ( TO_X01 ( DI1_ipd )    = 'X' ) or
          ( TO_X01 ( DI0_ipd )    = 'X' )
         ) then
        wpe_var  :=  'X';
      elsif ( TO_X01 ( WCLKS_ipd ) = '1' ) then
        if ( tmp_par2 /= PARODD_ipd ) then
          wpe_var  :=  '1';
        else
          wpe_var  :=  '0';
        end if;
      end if;
      RAM_di_int(8) := DI8_delayed;
      WPE_zd := wpe_var;
    end if;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

    if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
    end if; 

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

  if (TO_X01(WCLKS_ipd)='X') then
   if (TO_X01(WCLKS_previous) /= 'X') then
    assert false
    report ": WCLK unknown"
    severity Warning;
    end if;
   elsif (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      case TO_X01(WBint_delayed) is
          when '1' =>
            null;
          when '0' =>
           if(WADDR < 0) then
            if ((TO_X01(WADDR0_delayed) = 'X') and (TO_X01(WADDR0_previous) /= 'X')) then
             assert false
             report ": WADDR0 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR1_delayed) = 'X') and (TO_X01(WADDR1_previous) /= 'X')) then
             assert false
             report ": WADDR1 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR2_delayed) = 'X') and (TO_X01(WADDR2_previous) /= 'X')) then
             assert false
             report ": WADDR2 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR3_delayed) = 'X') and (TO_X01(WADDR3_previous) /= 'X')) then
             assert false
             report ": WADDR3 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR4_delayed) = 'X') and (TO_X01(WADDR4_previous) /= 'X')) then
             assert false
             report ": WADDR4 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR5_delayed) = 'X') and (TO_X01(WADDR5_previous) /= 'X')) then
             assert false
             report ": WADDR5 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR6_delayed) = 'X') and (TO_X01(WADDR6_previous) /= 'X')) then
             assert false
             report ": WADDR6 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR7_delayed) = 'X') and (TO_X01(WADDR7_previous) /= 'X')) then
             assert false
             report ": WADDR7 unknown"
             severity Warning;
            end if;
           else 
             RAM_di_int(7 downto 0) := DI7_delayed & DI6_delayed & DI5_delayed & DI4_delayed & DI3_delayed & DI2_delayed & DI1_delayed & DI0_delayed;
             memory_array(WADDR)  := RAM_di_int;
           end if;

         when others =>
          if (TO_X01(WBint_previous) /= 'X') then
             assert false
             report ": WRB or WBLKB unknown"
             severity Warning;
           end if;
      end case;
    end if;


 -----------------------------------------------------------
 --  Read Functional Section                              --
 -----------------------------------------------------------


    if (TO_X01(RCLKS_ipd) = 'X') then
       DO0_stg1 := 'X';
       DO1_stg1 := 'X';
       DO2_stg1 := 'X';
       DO3_stg1 := 'X';
       DO4_stg1 := 'X';
       DO5_stg1 := 'X';
       DO6_stg1 := 'X';
       DO7_stg1 := 'X';
       DO8_stg1 := 'X';
       RPE_stg1 := 'X';
       if (TO_X01(RCLKS_previous) /= 'X') then
         assert false
         report ": RCLK unknown"
         severity Warning;
       end if;
    elsif(RCLKS_ipd'event and RCLKS_ipd = '1') then

      DO0_zd := DO0_stg1;
      DO1_zd := DO1_stg1;
      DO2_zd := DO2_stg1;
      DO3_zd := DO3_stg1;
      DO4_zd := DO4_stg1;
      DO5_zd := DO5_stg1;
      DO6_zd := DO6_stg1;
      DO7_zd := DO7_stg1;
      DO8_zd := DO8_stg1;
      RPE_zd := RPE_stg1;

      case TO_X01(RBint_delayed) is
          when '1' =>
           null;
          when '0' =>

          if(RADDR < 0) then 
          DO0_stg1 := 'X';
          DO1_stg1 := 'X';
          DO2_stg1 := 'X';
          DO3_stg1 := 'X';
          DO4_stg1 := 'X';
          DO5_stg1 := 'X';
          DO6_stg1 := 'X';
          DO7_stg1 := 'X';
          DO8_stg1 := 'X';
          RPE_stg1 := 'X';
          if(TO_X01(RADDR0_delayed) = 'X') and (TO_X01(RADDR0_previous) /= 'X') then
             assert false
             report ": RADDR0 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR1_delayed) = 'X') and (TO_X01(RADDR1_previous) /= 'X') then
             assert false
             report ": RADDR1 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR2_delayed) = 'X') and (TO_X01(RADDR2_previous) /= 'X') then
             assert false
             report ": RADDR2 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR3_delayed) = 'X') and (TO_X01(RADDR3_previous) /= 'X') then
             assert false
             report ": RADDR3 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR4_delayed) = 'X') and (TO_X01(RADDR4_previous) /= 'X') then
             assert false
             report ": RADDR4 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR5_delayed) = 'X') and (TO_X01(RADDR5_previous) /= 'X') then
             assert false
             report ": RADDR5 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR6_delayed) = 'X') and (TO_X01(RADDR6_previous) /= 'X') then
             assert false
             report ": RADDR6 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR7_delayed) = 'X') and (TO_X01(RADDR7_previous) /= 'X') then
             assert false
             report ": RADDR7 unknown"
             severity Warning;
          end if;
          else  
            DO0_stg1 :=memory_array(RADDR)(0);
            DO1_stg1 :=memory_array(RADDR)(1);
            DO2_stg1 :=memory_array(RADDR)(2);
            DO3_stg1 :=memory_array(RADDR)(3);
            DO4_stg1 :=memory_array(RADDR)(4);
            DO5_stg1 :=memory_array(RADDR)(5);
            DO6_stg1 :=memory_array(RADDR)(6);
            DO7_stg1 :=memory_array(RADDR)(7);
            DO8_stg1 :=memory_array(RADDR)(8);
            do_par  := DO8_stg1 XOR DO7_stg1 XOR DO6_stg1 XOR DO5_stg1 XOR DO4_stg1 XOR DO3_stg1 XOR DO2_stg1 XOR DO1_stg1 XOR DO0_stg1;
            par_f <= do_par;
            if ( do_par = 'X' ) then
              RPE_stg1 := 'X';
            elsif ( TO_X01 ( PARODD_delayed ) = 'X' ) then
              RPE_stg1 := 'X';
            else
              if ( do_par /= PARODD_delayed ) then
                RPE_stg1  :=  '1';
              else
                RPE_stg1  :=  '0';
              end if;
            end if;
        end if;

         when others =>
          DO0_stg1 := 'X';
          DO1_stg1 := 'X';
          DO2_stg1 := 'X';
          DO3_stg1 := 'X';
          DO4_stg1 := 'X';
          DO5_stg1 := 'X';
          DO6_stg1 := 'X';
          DO7_stg1 := 'X';
          DO8_stg1 := 'X';
          RPE_stg1 := 'X';
          if(TO_X01(RBint_previous) /= 'X') then
             assert false
             report ": RDB or RBLKB unknown "
             severity Warning;
           end if;
         end case;
       end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       WCLKS_previous  := WCLKS_ipd;
       RCLKS_previous  := RCLKS_ipd;
       RBint_previous := RBint_delayed;
       RBint_delayed  := RBint;
       WBint_previous  := WBint_delayed;
       WBint_delayed   := WBint;
       DI0_delayed     := DI0_ipd;
       DI1_delayed     := DI1_ipd;
       DI2_delayed     := DI2_ipd;
       DI3_delayed     := DI3_ipd;
       DI4_delayed     := DI4_ipd;
       DI5_delayed     := DI5_ipd;
       DI6_delayed     := DI6_ipd;
       DI7_delayed     := DI7_ipd;
       DI8_delayed     := DI8_ipd;
       RADDR0_previous := RADDR0_delayed;
       RADDR0_delayed  := RADDR0_ipd;
       RADDR1_previous := RADDR1_delayed;
       RADDR1_delayed  := RADDR1_ipd;
       RADDR2_previous := RADDR2_delayed;
       RADDR2_delayed  := RADDR2_ipd;
       RADDR3_previous := RADDR3_delayed;
       RADDR3_delayed  := RADDR3_ipd;
       RADDR4_previous := RADDR4_delayed;
       RADDR4_delayed  := RADDR4_ipd;
       RADDR5_previous := RADDR5_delayed;
       RADDR5_delayed  := RADDR5_ipd;
       RADDR6_previous := RADDR6_delayed;
       RADDR6_delayed  := RADDR6_ipd;
       RADDR7_previous := RADDR7_delayed;
       RADDR7_delayed  := RADDR7_ipd;
       WADDR0_previous := WADDR0_delayed;
       WADDR0_delayed  := WADDR0_ipd;
       WADDR1_previous := WADDR1_delayed;
       WADDR1_delayed  := WADDR1_ipd;
       WADDR2_previous := WADDR2_delayed;
       WADDR2_delayed  := WADDR2_ipd;
       WADDR3_previous := WADDR3_delayed;
       WADDR3_delayed  := WADDR3_ipd;
       WADDR4_previous := WADDR4_delayed;
       WADDR4_delayed  := WADDR4_ipd;
       WADDR5_previous := WADDR5_delayed;
       WADDR5_delayed  := WADDR5_ipd;
       WADDR6_previous := WADDR6_delayed;
       WADDR6_delayed  := WADDR6_ipd;
       WADDR7_previous := WADDR7_delayed;
       WADDR7_delayed  := WADDR7_ipd;
       PARODD_previous := PARODD_delayed; 
       PARODD_delayed  := PARODD_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
           OutSignal     => DOS,
           GlitchData    => DOS_GlitchData,
           OutSignalName => "DOS",
           OutTemp       => DOS_zd,
           Paths  =>  (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),
           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
             OutSignal     => WPE,
             GlitchData    => WPE_GlitchData,
             OutSignalName => "WPE",
             OutTemp       => WPE_zd,
             Paths =>   (0 => (WCLKS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_WCLKS_WPE), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
         OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => RPE,
           GlitchData    => RPE_GlitchData,
           OutSignalName => "RPE",
           OutTemp       => RPE_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_RPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
LIBRARY STD;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

USE std.textio.all;
USE ieee.std_logic_textio.all;
LIBRARY a500k;
USE a500k.all;

entity RAM256x9SSRP is 

   generic (
        Xon                     : Boolean := False;
        MsgOn                   : Boolean := True;
        TimingCheckOn           : Boolean := True;
        MEMORYFILE              : String  := "";
        InstancePath            : String  := "*";

 	tipd_RADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WADDR7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tsetup_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RDB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR0_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR0_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR1_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR1_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR2_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR2_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR3_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR3_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR4_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR4_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR5_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR5_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR6_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR6_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RADDR7_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RADDR7_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge	                : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge	                : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS	                        : VitalDelayType := 0.000 ns;
 	tsetup_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR0_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR0_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR1_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR1_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR2_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR2_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR3_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR3_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR4_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR4_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR5_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR5_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR6_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR6_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WADDR7_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WADDR7_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_negedge_posedge	        : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_posedge_posedge	        : VitalDelayType := 0.000 ns;
	tpw_WCLKS_posedge                       : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                       : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                           : VitalDelayType := 0.000 ns;

 	-- timing data for checking read/write at the same address, and at same time
 	tsetup_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 0.000 ns;
 	thold_WCLKS_RCLKS_posedge_posedge	: VitalDelayType := 7.000 ns

 	);
 port (
   DO0    :  OUT STD_LOGIC := 'X';
   DO1    :  OUT STD_LOGIC := 'X';
   DO2    :  OUT STD_LOGIC := 'X';
   DO3    :  OUT STD_LOGIC := 'X';
   DO4    :  OUT STD_LOGIC := 'X';
   DO5    :  OUT STD_LOGIC := 'X';
   DO6    :  OUT STD_LOGIC := 'X';
   DO7    :  OUT STD_LOGIC := 'X';
   DO8    :  OUT STD_LOGIC := 'X';
   DOS    :  OUT STD_LOGIC := 'X';

   WADDR0 :  IN STD_LOGIC := 'X';
   WADDR1 :  IN STD_LOGIC := 'X';
   WADDR2 :  IN STD_LOGIC := 'X';
   WADDR3 :  IN STD_LOGIC := 'X';
   WADDR4 :  IN STD_LOGIC := 'X';
   WADDR5 :  IN STD_LOGIC := 'X';
   WADDR6 :  IN STD_LOGIC := 'X';
   WADDR7 :  IN STD_LOGIC := 'X';
   RADDR0 :  IN STD_LOGIC := 'X';
   RADDR1 :  IN STD_LOGIC := 'X';
   RADDR2 :  IN STD_LOGIC := 'X';
   RADDR3 :  IN STD_LOGIC := 'X';
   RADDR4 :  IN STD_LOGIC := 'X';
   RADDR5 :  IN STD_LOGIC := 'X';
   RADDR6 :  IN STD_LOGIC := 'X';
   RADDR7 :  IN STD_LOGIC := 'X';
   DI0    :  IN STD_LOGIC := 'X';
   DI1    :  IN STD_LOGIC := 'X';
   DI2    :  IN STD_LOGIC := 'X';
   DI3    :  IN STD_LOGIC := 'X';
   DI4    :  IN STD_LOGIC := 'X';
   DI5    :  IN STD_LOGIC := 'X';
   DI6    :  IN STD_LOGIC := 'X';
   DI7    :  IN STD_LOGIC := 'X';
   DI8    :  IN STD_LOGIC := 'X';
   WRB    :  IN STD_LOGIC := 'X';
   RDB    :  IN STD_LOGIC := 'X';
   WBLKB  :  IN STD_LOGIC := 'X';
   RBLKB  :  IN STD_LOGIC := 'X';
   PARODD :  IN STD_LOGIC := 'X';
   RCLKS   :  IN STD_LOGIC := 'X';
   WCLKS   :  IN STD_LOGIC := 'X';
   DIS    :  IN STD_LOGIC := 'X');

ATTRIBUTE VITAL_LEVEL0 OF RAM256x9SSRP : entity IS True ;
END RAM256x9SSRP;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of RAM256x9SSRP is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal WADDR0_ipd : std_ulogic := 'X';
   signal WADDR1_ipd : std_ulogic := 'X';
   signal WADDR2_ipd : std_ulogic := 'X';
   signal WADDR3_ipd : std_ulogic := 'X';
   signal WADDR4_ipd : std_ulogic := 'X';
   signal WADDR5_ipd : std_ulogic := 'X';
   signal WADDR6_ipd : std_ulogic := 'X';
   signal WADDR7_ipd : std_ulogic := 'X';
   signal RADDR0_ipd : std_ulogic := 'X';
   signal RADDR1_ipd : std_ulogic := 'X';
   signal RADDR2_ipd : std_ulogic := 'X';
   signal RADDR3_ipd : std_ulogic := 'X';
   signal RADDR4_ipd : std_ulogic := 'X';
   signal RADDR5_ipd : std_ulogic := 'X';
   signal RADDR6_ipd : std_ulogic := 'X';
   signal RADDR7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal WCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

	-- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';
   signal INIT_MEM   : std_logic:= '0';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic:= 'X';
   signal par_f2     : std_logic:= 'X';

 begin  --  VITAL_ACT
   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (WADDR0_ipd, WADDR0, VitalExtendToFillDelay(tipd_WADDR0));
   VitalWireDelay (WADDR1_ipd, WADDR1, VitalExtendToFillDelay(tipd_WADDR1));
   VitalWireDelay (WADDR2_ipd, WADDR2, VitalExtendToFillDelay(tipd_WADDR2));
   VitalWireDelay (WADDR3_ipd, WADDR3, VitalExtendToFillDelay(tipd_WADDR3));
   VitalWireDelay (WADDR4_ipd, WADDR4, VitalExtendToFillDelay(tipd_WADDR4));
   VitalWireDelay (WADDR5_ipd, WADDR5, VitalExtendToFillDelay(tipd_WADDR5));
   VitalWireDelay (WADDR6_ipd, WADDR6, VitalExtendToFillDelay(tipd_WADDR6));
   VitalWireDelay (WADDR7_ipd, WADDR7, VitalExtendToFillDelay(tipd_WADDR7));
   VitalWireDelay (RADDR0_ipd, RADDR0, VitalExtendToFillDelay(tipd_RADDR0));
   VitalWireDelay (RADDR1_ipd, RADDR1, VitalExtendToFillDelay(tipd_RADDR1));
   VitalWireDelay (RADDR2_ipd, RADDR2, VitalExtendToFillDelay(tipd_RADDR2));
   VitalWireDelay (RADDR3_ipd, RADDR3, VitalExtendToFillDelay(tipd_RADDR3));
   VitalWireDelay (RADDR4_ipd, RADDR4, VitalExtendToFillDelay(tipd_RADDR4));
   VitalWireDelay (RADDR5_ipd, RADDR5, VitalExtendToFillDelay(tipd_RADDR5));
   VitalWireDelay (RADDR6_ipd, RADDR6, VitalExtendToFillDelay(tipd_RADDR6));
   VitalWireDelay (RADDR7_ipd, RADDR7, VitalExtendToFillDelay(tipd_RADDR7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (WCLKS_ipd, WCLKS, VitalExtendToFillDelay(tipd_WCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

---------------------------------------------------------------
--                  Behavior Section                         --
---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);


    PROCESS
    BEGIN
      INIT_MEM <= '1';
      WAIT;
    END PROCESS;

    VITALBehavior : process (INIT_MEM, 
                          RADDR0_ipd, RADDR1_ipd, RADDR2_ipd, RADDR3_ipd, RADDR4_ipd, RADDR5_ipd, RADDR6_ipd, RADDR7_ipd, 
                          WADDR0_ipd, WADDR1_ipd, WADDR2_ipd, WADDR3_ipd, WADDR4_ipd, WADDR5_ipd, WADDR6_ipd, WADDR7_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd 
                          )

    -- some internal veriable declaration
     variable RAM_di_int         : std_logic_vector(8 downto 0);
     variable memory_array       : MEM_TYPE := (others =>(others => 'X'));
     variable do_par             : std_logic:= 'X';
     variable tmp_par            : std_logic:= 'X';
     variable tmp_par2           : std_logic:= 'X';
     variable wpe_var            : std_logic:= 'X';

     --  Read Timing Check Results
     variable Tviol_RADDR0_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR0_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR1_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR1_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR2_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR2_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR3_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR3_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR4_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR4_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR5_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR5_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR6_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR6_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RADDR7_RCLKS_posedge : X01                 := '0';
     variable TmDt_RADDR7_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable Tviol_WADDR0_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR0_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR1_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR1_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR2_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR2_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR3_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR3_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR4_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR4_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR5_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR5_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR6_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR6_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WADDR7_WCLKS_posedge : X01                 := '0';
     variable TmDt_WADDR7_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI0_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI1_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI2_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI3_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI4_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI5_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI6_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI7_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI8_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_WCLKS_posedge    : X01                 := '0';
     variable TmDt_WRB_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_WCLKS_posedge  : X01                 := '0';
     variable TmDt_WBLKB_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WCLKS                : X01                 := '0';
     variable Tviol_WCLKS_RCLKS_posedge  : X01                 := '0';
     variable TmDt_WCLKS_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results

     variable WADDR : integer := -1;
     variable RADDR : integer := -1;
     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     variable DO0_zd : std_ulogic;
     variable DO1_zd : std_ulogic;
     variable DO2_zd : std_ulogic;
     variable DO3_zd : std_ulogic;
     variable DO4_zd : std_ulogic;
     variable DO5_zd : std_ulogic;
     variable DO6_zd : std_ulogic;
     variable DO7_zd : std_ulogic;
     variable DO8_zd : std_ulogic;
     variable RPE_zd : std_ulogic;
     variable WPE_zd : std_ulogic;
     variable DOS_zd : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData  : VitalGlitchDataType;
     variable DO1_GlitchData  : VitalGlitchDataType;
     variable DO2_GlitchData  : VitalGlitchDataType;
     variable DO3_GlitchData  : VitalGlitchDataType;
     variable DO4_GlitchData  : VitalGlitchDataType;
     variable DO5_GlitchData  : VitalGlitchDataType;
     variable DO6_GlitchData  : VitalGlitchDataType;
     variable DO7_GlitchData  : VitalGlitchDataType;
     variable DO8_GlitchData  : VitalGlitchDataType;
     variable DOS_GlitchData  : VitalGlitchDataType;

     -- last value variables
     variable WCLKS_previous  : std_ulogic := 'X';
     variable RCLKS_previous  : std_ulogic := 'X';
     variable RBint_delayed   : std_ulogic := 'X';
     variable RBint_previous  : std_ulogic := 'X';
     variable WBint_delayed   : std_ulogic := 'X';
     variable WBint_previous  : std_ulogic := 'X';
     variable DIS_previous    : std_ulogic := 'X';
     variable DI0_delayed     : std_ulogic := 'X';
     variable DI1_delayed     : std_ulogic := 'X';
     variable DI2_delayed     : std_ulogic := 'X';
     variable DI3_delayed     : std_ulogic := 'X';
     variable DI4_delayed     : std_ulogic := 'X';
     variable DI5_delayed     : std_ulogic := 'X';
     variable DI6_delayed     : std_ulogic := 'X';
     variable DI7_delayed     : std_ulogic := 'X';
     variable DI8_delayed     : std_ulogic := 'X';
     variable RADDR0_delayed  : std_ulogic := 'X';
     variable RADDR1_delayed  : std_ulogic := 'X';
     variable RADDR2_delayed  : std_ulogic := 'X';
     variable RADDR3_delayed  : std_ulogic := 'X';
     variable RADDR4_delayed  : std_ulogic := 'X';
     variable RADDR5_delayed  : std_ulogic := 'X';
     variable RADDR6_delayed  : std_ulogic := 'X';
     variable RADDR7_delayed  : std_ulogic := 'X';
     variable RADDR0_previous : std_ulogic := 'X';
     variable RADDR1_previous : std_ulogic := 'X';
     variable RADDR2_previous : std_ulogic := 'X';
     variable RADDR3_previous : std_ulogic := 'X';
     variable RADDR4_previous : std_ulogic := 'X';
     variable RADDR5_previous : std_ulogic := 'X';
     variable RADDR6_previous : std_ulogic := 'X';
     variable RADDR7_previous : std_ulogic := 'X';
     variable WADDR0_delayed  : std_ulogic := 'X';
     variable WADDR1_delayed  : std_ulogic := 'X';
     variable WADDR2_delayed  : std_ulogic := 'X';
     variable WADDR3_delayed  : std_ulogic := 'X';
     variable WADDR4_delayed  : std_ulogic := 'X';
     variable WADDR5_delayed  : std_ulogic := 'X';
     variable WADDR6_delayed  : std_ulogic := 'X';
     variable WADDR7_delayed  : std_ulogic := 'X';
     variable WADDR0_previous : std_ulogic := 'X';
     variable WADDR1_previous : std_ulogic := 'X';
     variable WADDR2_previous : std_ulogic := 'X';
     variable WADDR3_previous : std_ulogic := 'X';
     variable WADDR4_previous : std_ulogic := 'X';
     variable WADDR5_previous : std_ulogic := 'X';
     variable WADDR6_previous : std_ulogic := 'X';
     variable WADDR7_previous : std_ulogic := 'X';

     --  Pipelined temporary results
     variable RPE_stg1        : std_ulogic := 'X';
     variable DO0_stg1        : std_ulogic := 'X';
     variable DO1_stg1        : std_ulogic := 'X';
     variable DO2_stg1        : std_ulogic := 'X';
     variable DO3_stg1        : std_ulogic := 'X';
     variable DO4_stg1        : std_ulogic := 'X';
     variable DO5_stg1        : std_ulogic := 'X';
     variable DO6_stg1        : std_ulogic := 'X';
     variable DO7_stg1        : std_ulogic := 'X';
     variable DO8_stg1        : std_ulogic := 'X';

     variable PARODD_delayed  : std_ulogic := 'X';
     variable PARODD_previous : std_ulogic := 'X';

     variable inline    : LINE;
     variable indata    : std_logic_vector(8 downto 0);
     variable resdata   : std_logic_vector(8 downto 0);
     variable i         : integer:=0;
     file     memfile   : text;
     variable status         : file_open_status;

 begin -- process VITALBehavior

  -----------------------------------------------------------
  --    Initialize memory file from MEMORYFILE string      --
  -----------------------------------------------------------


  if ( INIT_MEM'EVENT and INIT_MEM = '1') then
    file_open(status, memfile, MEMORYFILE, read_mode);
    if ( status=open_ok ) then
      while((i < 256) and (not ENDFILE(memfile))) loop
        readline(memfile,inline);
        read(inline,indata);
        resdata := indata;
        memory_array(i) := resdata;
        i := i+1;
      end loop;
    else
      assert ( MEMORYFILE'length = 0 )
        report "Failed to open RAM256x9SSRP memory initialization file in read mode"
        severity Note;
    end if;
    file_close(memfile);
  end if;

     if (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      WADDR := ((INT(WADDR7_delayed)*128)+(INT(WADDR6_delayed)*64)+(INT(
               WADDR5_delayed)*32) + (INT(WADDR4_delayed)*16) + 
               (INT(WADDR3_delayed)*8) + (INT(WADDR2_delayed)*4) + (INT(
               WADDR1_delayed)*2) + (INT(WADDR0_delayed)*1));
     end if;

   -- Convert Read Address Signal to Integer
     if (RCLKS_ipd'EVENT AND RCLKS_ipd = '1') then
      RADDR := ((INT(RADDR7_delayed)*128)+(INT(RADDR6_delayed)*64)+(INT(
               RADDR5_delayed)*32) + (INT(RADDR4_delayed)*16) + 
               (INT(RADDR3_delayed)*8) + (INT(RADDR2_delayed)*4) + (INT(
               RADDR1_delayed)*2) + (INT(RADDR0_delayed)*1));
     end if;

if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             tsetup_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             thold_RADDR0_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR0_RCLKS_posedge,
                             TmDt_RADDR0_RCLKS_posedge,
                             RADDR0_ipd, "RADDR0",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             tsetup_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             thold_RADDR0_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             tsetup_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             thold_RADDR1_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR1_RCLKS_posedge,
                             TmDt_RADDR1_RCLKS_posedge,
                             RADDR1_ipd, "RADDR1",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             tsetup_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             thold_RADDR1_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             tsetup_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             thold_RADDR2_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR2_RCLKS_posedge,
                             TmDt_RADDR2_RCLKS_posedge,
                             RADDR2_ipd, "RADDR2",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             tsetup_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             thold_RADDR2_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             tsetup_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             thold_RADDR3_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR3_RCLKS_posedge,
                             TmDt_RADDR3_RCLKS_posedge,
                             RADDR3_ipd, "RADDR3",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             tsetup_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             thold_RADDR3_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             tsetup_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             thold_RADDR4_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR4_RCLKS_posedge,
                             TmDt_RADDR4_RCLKS_posedge,
                             RADDR4_ipd, "RADDR4",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             tsetup_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             thold_RADDR4_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             tsetup_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             thold_RADDR5_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR5_RCLKS_posedge,
                             TmDt_RADDR5_RCLKS_posedge,
                             RADDR5_ipd, "RADDR5",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             tsetup_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             thold_RADDR5_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             tsetup_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             thold_RADDR6_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR6_RCLKS_posedge,
                             TmDt_RADDR6_RCLKS_posedge,
                             RADDR6_ipd, "RADDR6",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             tsetup_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             thold_RADDR6_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             tsetup_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             thold_RADDR7_RCLKS_posedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RADDR7_RCLKS_posedge,
                             TmDt_RADDR7_RCLKS_posedge,
                             RADDR7_ipd, "RADDR7",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             tsetup_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             thold_RADDR7_RCLKS_negedge_posedge,
                             (To_X01(RBint) = '0'),
                             '/',
                             InstancePath &" /RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

 -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             (To_X01(RBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             (To_X01(RDB_ipd) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (To_X01(RBLKB_ipd) = '0') AND (To_X01(RDB_ipd) = '0'),
                             InstancePath & "/RAM256x9SSRP",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       VitalSetupHoldCheck ( Tviol_WADDR0_WCLKS_posedge,
                             TmDt_WADDR0_WCLKS_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR0_WCLKS_posedge_posedge,
                             tsetup_WADDR0_WCLKS_posedge_posedge,
                             thold_WADDR0_WCLKS_posedge_posedge,
                             thold_WADDR0_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR0_WCLKS_posedge,
                             TmDt_WADDR0_WCLKS_posedge,
                             WADDR0_ipd, "WADDR0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR0_WCLKS_negedge_posedge,
                             tsetup_WADDR0_WCLKS_negedge_posedge,
                             thold_WADDR0_WCLKS_negedge_posedge,
                             thold_WADDR0_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WCLKS_posedge,
                             TmDt_WADDR1_WCLKS_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR1_WCLKS_posedge_posedge,
                             tsetup_WADDR1_WCLKS_posedge_posedge,
                             thold_WADDR1_WCLKS_posedge_posedge,
                             thold_WADDR1_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR1_WCLKS_posedge,
                             TmDt_WADDR1_WCLKS_posedge,
                             WADDR1_ipd, "WADDR1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR1_WCLKS_negedge_posedge,
                             tsetup_WADDR1_WCLKS_negedge_posedge,
                             thold_WADDR1_WCLKS_negedge_posedge,
                             thold_WADDR1_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WCLKS_posedge,
                             TmDt_WADDR2_WCLKS_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR2_WCLKS_posedge_posedge,
                             tsetup_WADDR2_WCLKS_posedge_posedge,
                             thold_WADDR2_WCLKS_posedge_posedge,
                             thold_WADDR2_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR2_WCLKS_posedge,
                             TmDt_WADDR2_WCLKS_posedge,
                             WADDR2_ipd, "WADDR2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR2_WCLKS_negedge_posedge,
                             tsetup_WADDR2_WCLKS_negedge_posedge,
                             thold_WADDR2_WCLKS_negedge_posedge,
                             thold_WADDR2_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WCLKS_posedge,
                             TmDt_WADDR3_WCLKS_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR3_WCLKS_posedge_posedge,
                             tsetup_WADDR3_WCLKS_posedge_posedge,
                             thold_WADDR3_WCLKS_posedge_posedge,
                             thold_WADDR3_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR3_WCLKS_posedge,
                             TmDt_WADDR3_WCLKS_posedge,
                             WADDR3_ipd, "WADDR3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR3_WCLKS_negedge_posedge,
                             tsetup_WADDR3_WCLKS_negedge_posedge,
                             thold_WADDR3_WCLKS_negedge_posedge,
                             thold_WADDR3_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WCLKS_posedge,
                             TmDt_WADDR4_WCLKS_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR4_WCLKS_posedge_posedge,
                             tsetup_WADDR4_WCLKS_posedge_posedge,
                             thold_WADDR4_WCLKS_posedge_posedge,
                             thold_WADDR4_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR4_WCLKS_posedge,
                             TmDt_WADDR4_WCLKS_posedge,
                             WADDR4_ipd, "WADDR4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR4_WCLKS_negedge_posedge,
                             tsetup_WADDR4_WCLKS_negedge_posedge,
                             thold_WADDR4_WCLKS_negedge_posedge,
                             thold_WADDR4_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WCLKS_posedge,
                             TmDt_WADDR5_WCLKS_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR5_WCLKS_posedge_posedge,
                             tsetup_WADDR5_WCLKS_posedge_posedge,
                             thold_WADDR5_WCLKS_posedge_posedge,
                             thold_WADDR5_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR5_WCLKS_posedge,
                             TmDt_WADDR5_WCLKS_posedge,
                             WADDR5_ipd, "WADDR5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR5_WCLKS_negedge_posedge,
                             tsetup_WADDR5_WCLKS_negedge_posedge,
                             thold_WADDR5_WCLKS_negedge_posedge,
                             thold_WADDR5_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WCLKS_posedge,
                             TmDt_WADDR6_WCLKS_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR6_WCLKS_posedge_posedge,
                             tsetup_WADDR6_WCLKS_posedge_posedge,
                             thold_WADDR6_WCLKS_posedge_posedge,
                             thold_WADDR6_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR6_WCLKS_posedge,
                             TmDt_WADDR6_WCLKS_posedge,
                             WADDR6_ipd, "WADDR6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR6_WCLKS_negedge_posedge,
                             tsetup_WADDR6_WCLKS_negedge_posedge,
                             thold_WADDR6_WCLKS_negedge_posedge,
                             thold_WADDR6_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WCLKS_posedge,
                             TmDt_WADDR7_WCLKS_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR7_WCLKS_posedge_posedge,
                             tsetup_WADDR7_WCLKS_posedge_posedge,
                             thold_WADDR7_WCLKS_posedge_posedge,
                             thold_WADDR7_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WADDR7_WCLKS_posedge,
                             TmDt_WADDR7_WCLKS_posedge,
                             WADDR7_ipd, "WADDR7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WADDR7_WCLKS_negedge_posedge,
                             tsetup_WADDR7_WCLKS_negedge_posedge,
                             thold_WADDR7_WCLKS_negedge_posedge,
                             thold_WADDR7_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath &"/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_posedge_posedge,
                             tsetup_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_negedge_posedge,
                             tsetup_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_posedge_posedge,
                             tsetup_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_negedge_posedge,
                             tsetup_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_posedge_posedge,
                             tsetup_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_negedge_posedge,
                             tsetup_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_posedge_posedge,
                             tsetup_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_negedge_posedge,
                             tsetup_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_posedge_posedge,
                             tsetup_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_negedge_posedge,
                             tsetup_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_posedge_posedge,
                             tsetup_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_negedge_posedge,
                             tsetup_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_posedge_posedge,
                             tsetup_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_negedge_posedge,
                             tsetup_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_posedge_posedge,
                             tsetup_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_negedge_posedge,
                             tsetup_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_posedge_posedge,
                             tsetup_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_negedge_posedge,
                             tsetup_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             (To_X01(WBint) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

 -- setup hold WEN, WBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_posedge_posedge,
                             tsetup_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_negedge_posedge,
                             tsetup_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             (To_X01(WBLKB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             (To_X01(WRB_ipd) = '0'),
                             '/',
                             InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

  --   Period of WCLK
      VitalPeriodPulseCheck ( Pviol_WCLKS,
                              PeriodData_WCLKS,
                              WCLKS_ipd, "WCLKS",
                              0.0 ns,
                              tperiod_WCLKS,
                              tpw_WCLKS_posedge,
                              tpw_WCLKS_negedge,
                              (To_X01(WBLKB_ipd) = '0') AND (To_X01(WRB_ipd) = '0'),
                             InstancePath & "/RAM256x9SSRP",
                              True,
                              True,
                              WARNING
                              );
   ------------------------------------------------------------
   --        Timing Checking for Read and write conflict     --
   ------------------------------------------------------------
       VitalSetupHoldCheck ( Tviol_WCLKS_RCLKS_posedge,
                             TmDt_WCLKS_RCLKS_posedge,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_WCLKS_RCLKS_posedge_posedge,
                             0.0 ns,
                             thold_WCLKS_RCLKS_posedge_posedge,
                             0.0 ns,
                             (To_X01(RBint) = '0') AND (To_X01(WBint) = '0') AND (RADDR = WADDR),
                             '/',
                              InstancePath & "/RAM256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

 end if;

   ------------------------------------------------------------
   --         WPE generating  block                            -
   ------------------------------------------------------------

     if (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
        tmp_par  := DI7_delayed XOR DI6_delayed XOR DI5_delayed XOR DI4_delayed XOR DI3_delayed XOR DI2_delayed XOR DI1_delayed XOR DI0_delayed;
        if (tmp_par   /= PARODD_delayed) then
           wpe_var     :=  '1';
        else
           wpe_var     :=  '0';
        end if;
        RAM_di_int(8) := wpe_var;
        WPE_zd := wpe_var;
     end if;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

    if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
    end if; 

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

  if (TO_X01(WCLKS_ipd)='X') then
   if (TO_X01(WCLKS_previous) /= 'X') then
    assert false
    report ": WCLK unknown"
    severity Warning;
    end if;
   elsif (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      case TO_X01(WBint_delayed) is
          when '1' =>
            null;
          when '0' =>
           if(WADDR < 0) then
            if ((TO_X01(WADDR0_delayed) = 'X') and (TO_X01(WADDR0_previous) /= 'X')) then
             assert false
             report ": WADDR0 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR1_delayed) = 'X') and (TO_X01(WADDR1_previous) /= 'X')) then
             assert false
             report ": WADDR1 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR2_delayed) = 'X') and (TO_X01(WADDR2_previous) /= 'X')) then
             assert false
             report ": WADDR2 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR3_delayed) = 'X') and (TO_X01(WADDR3_previous) /= 'X')) then
             assert false
             report ": WADDR3 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR4_delayed) = 'X') and (TO_X01(WADDR4_previous) /= 'X')) then
             assert false
             report ": WADDR4 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR5_delayed) = 'X') and (TO_X01(WADDR5_previous) /= 'X')) then
             assert false
             report ": WADDR5 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR6_delayed) = 'X') and (TO_X01(WADDR6_previous) /= 'X')) then
             assert false
             report ": WADDR6 unknown"
             severity Warning;
            end if;
            if ((TO_X01(WADDR7_delayed) = 'X') and (TO_X01(WADDR7_previous) /= 'X')) then
             assert false
             report ": WADDR7 unknown"
             severity Warning;
            end if;
           else 
             RAM_di_int(7 downto 0) := DI7_delayed & DI6_delayed & DI5_delayed & DI4_delayed & DI3_delayed & DI2_delayed & DI1_delayed & DI0_delayed;
             memory_array(WADDR)  := RAM_di_int;
           end if;

         when others =>
          if (TO_X01(WBint_previous) /= 'X') then
             assert false
             report ": WRB or WBLKB unknown"
             severity Warning;
           end if;
      end case;
    end if;


 -----------------------------------------------------------
 --  Read Functional Section                              --
 -----------------------------------------------------------


    if (TO_X01(RCLKS_ipd) = 'X') then
       DO0_stg1 := 'X';
       DO1_stg1 := 'X';
       DO2_stg1 := 'X';
       DO3_stg1 := 'X';
       DO4_stg1 := 'X';
       DO5_stg1 := 'X';
       DO6_stg1 := 'X';
       DO7_stg1 := 'X';
       DO8_stg1 := 'X';
       RPE_stg1 := 'X';
       if (TO_X01(RCLKS_previous) /= 'X') then
         assert false
         report ": RCLK unknown"
         severity Warning;
       end if;
    elsif(RCLKS_ipd'event and RCLKS_ipd = '1') then

      DO0_zd := DO0_stg1;
      DO1_zd := DO1_stg1;
      DO2_zd := DO2_stg1;
      DO3_zd := DO3_stg1;
      DO4_zd := DO4_stg1;
      DO5_zd := DO5_stg1;
      DO6_zd := DO6_stg1;
      DO7_zd := DO7_stg1;
      DO8_zd := DO8_stg1;
      RPE_zd := RPE_stg1;

      case TO_X01(RBint_delayed) is
          when '1' =>
           null;
          when '0' =>

          if(RADDR < 0) then 
          DO0_stg1 := 'X';
          DO1_stg1 := 'X';
          DO2_stg1 := 'X';
          DO3_stg1 := 'X';
          DO4_stg1 := 'X';
          DO5_stg1 := 'X';
          DO6_stg1 := 'X';
          DO7_stg1 := 'X';
          DO8_stg1 := 'X';
          if(TO_X01(RADDR0_delayed) = 'X') and (TO_X01(RADDR0_previous) /= 'X') then
             assert false
             report ": RADDR0 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR1_delayed) = 'X') and (TO_X01(RADDR1_previous) /= 'X') then
             assert false
             report ": RADDR1 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR2_delayed) = 'X') and (TO_X01(RADDR2_previous) /= 'X') then
             assert false
             report ": RADDR2 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR3_delayed) = 'X') and (TO_X01(RADDR3_previous) /= 'X') then
             assert false
             report ": RADDR3 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR4_delayed) = 'X') and (TO_X01(RADDR4_previous) /= 'X') then
             assert false
             report ": RADDR4 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR5_delayed) = 'X') and (TO_X01(RADDR5_previous) /= 'X') then
             assert false
             report ": RADDR5 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR6_delayed) = 'X') and (TO_X01(RADDR6_previous) /= 'X') then
             assert false
             report ": RADDR6 unknown"
             severity Warning;
          end if;
          if(TO_X01(RADDR7_delayed) = 'X') and (TO_X01(RADDR7_previous) /= 'X') then
             assert false
             report ": RADDR7 unknown"
             severity Warning;
          end if;
          else  
            DO0_stg1 :=memory_array(RADDR)(0);
            DO1_stg1 :=memory_array(RADDR)(1);
            DO2_stg1 :=memory_array(RADDR)(2);
            DO3_stg1 :=memory_array(RADDR)(3);
            DO4_stg1 :=memory_array(RADDR)(4);
            DO5_stg1 :=memory_array(RADDR)(5);
            DO6_stg1 :=memory_array(RADDR)(6);
            DO7_stg1 :=memory_array(RADDR)(7);
            DO8_stg1 :=memory_array(RADDR)(8);
        end if;

         when others =>
          DO0_stg1 := 'X';
          DO1_stg1 := 'X';
          DO2_stg1 := 'X';
          DO3_stg1 := 'X';
          DO4_stg1 := 'X';
          DO5_stg1 := 'X';
          DO6_stg1 := 'X';
          DO7_stg1 := 'X';
          DO8_stg1 := 'X';
          if(TO_X01(RBint_previous) /= 'X') then
             assert false
             report ": RDB or RBLKB unknown "
             severity Warning;
           end if;
         end case;
       end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       WCLKS_previous  := WCLKS_ipd;
       RCLKS_previous  := RCLKS_ipd;
       RBint_previous := RBint_delayed;
       RBint_delayed  := RBint;
       WBint_previous  := WBint_delayed;
       WBint_delayed   := WBint;
       DI0_delayed     := DI0_ipd;
       DI1_delayed     := DI1_ipd;
       DI2_delayed     := DI2_ipd;
       DI3_delayed     := DI3_ipd;
       DI4_delayed     := DI4_ipd;
       DI5_delayed     := DI5_ipd;
       DI6_delayed     := DI6_ipd;
       DI7_delayed     := DI7_ipd;
       DI8_delayed     := DI8_ipd;
       RADDR0_previous := RADDR0_delayed;
       RADDR0_delayed  := RADDR0_ipd;
       RADDR1_previous := RADDR1_delayed;
       RADDR1_delayed  := RADDR1_ipd;
       RADDR2_previous := RADDR2_delayed;
       RADDR2_delayed  := RADDR2_ipd;
       RADDR3_previous := RADDR3_delayed;
       RADDR3_delayed  := RADDR3_ipd;
       RADDR4_previous := RADDR4_delayed;
       RADDR4_delayed  := RADDR4_ipd;
       RADDR5_previous := RADDR5_delayed;
       RADDR5_delayed  := RADDR5_ipd;
       RADDR6_previous := RADDR6_delayed;
       RADDR6_delayed  := RADDR6_ipd;
       RADDR7_previous := RADDR7_delayed;
       RADDR7_delayed  := RADDR7_ipd;
       WADDR0_previous := WADDR0_delayed;
       WADDR0_delayed  := WADDR0_ipd;
       WADDR1_previous := WADDR1_delayed;
       WADDR1_delayed  := WADDR1_ipd;
       WADDR2_previous := WADDR2_delayed;
       WADDR2_delayed  := WADDR2_ipd;
       WADDR3_previous := WADDR3_delayed;
       WADDR3_delayed  := WADDR3_ipd;
       WADDR4_previous := WADDR4_delayed;
       WADDR4_delayed  := WADDR4_ipd;
       WADDR5_previous := WADDR5_delayed;
       WADDR5_delayed  := WADDR5_ipd;
       WADDR6_previous := WADDR6_delayed;
       WADDR6_delayed  := WADDR6_ipd;
       WADDR7_previous := WADDR7_delayed;
       WADDR7_delayed  := WADDR7_ipd;
       PARODD_previous := PARODD_delayed; 
       PARODD_delayed  := PARODD_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
           OutSignal     => DOS,
           GlitchData    => DOS_GlitchData,
           OutSignalName => "DOS",
           OutTemp       => DOS_zd,
           Paths  =>  (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),
           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
         OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths  =>  (0 => (RCLKS_ipd'last_event,
                                 VitalExtendToFillDelay(tpd_RCLKS_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );


   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

LIBRARY a500k;
USE a500k.all;

entity FIFO256x9AA is 
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI0_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI1_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI2_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI3_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI4_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI5_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI6_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI7_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI8_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tpw_RDB_posedge         : VitalDelayType        := 0.000 ns;
 	tpw_RDB_negedge         : VitalDelayType        := 0.000 ns;
 	tperiod_RDB             : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_posedge       : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_negedge       : VitalDelayType        := 0.000 ns;
 	tperiod_RBLKB           : VitalDelayType        := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;

  	-- WB falling edge hold to RESETB   
 	thold_WRB_RESET_posedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_RESET_posedge_posedge             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_RESET_posedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RESET_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_WRB_RESET_negedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WBLKB_RESET_negedge_posedge             : VitalDelayType := 0.000 ns;
	tsetup_WRB_RESET_negedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_RESET_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                               : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                               : VitalDelayType := 0.000 ns;
 	tperiod_WRB                                   : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        WPE    :  OUT STD_LOGIC := 'X';
        RPE    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');


ATTRIBUTE VITAL_LEVEL0 OF FIFO256x9AA : entity IS True ;
END FIFO256x9AA;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of FIFO256x9AA is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal LGDEP0_ipd : std_ulogic := 'X';
   signal LGDEP1_ipd : std_ulogic := 'X';
   signal LGDEP2_ipd : std_ulogic := 'X';
   signal LEVEL0_ipd : std_ulogic := 'X';
   signal LEVEL1_ipd : std_ulogic := 'X';
   signal LEVEL2_ipd : std_ulogic := 'X';
   signal LEVEL3_ipd : std_ulogic := 'X';
   signal LEVEL4_ipd : std_ulogic := 'X';
   signal LEVEL5_ipd : std_ulogic := 'X';
   signal LEVEL6_ipd : std_ulogic := 'X';
   signal LEVEL7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal RESET_ipd  : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

   -- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic := 'X';
   signal par_f2     : std_logic := 'X';

   signal WRITE_AT_PREV_EDGE : std_logic := '0';
   signal READ_AT_PREV_EDGE  : std_logic := '0';
   

   begin  --  VITAL_ACT

   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (LGDEP0_ipd, LGDEP0, VitalExtendToFillDelay(tipd_LGDEP0));
   VitalWireDelay (LGDEP1_ipd, LGDEP1, VitalExtendToFillDelay(tipd_LGDEP1));
   VitalWireDelay (LGDEP2_ipd, LGDEP2, VitalExtendToFillDelay(tipd_LGDEP2));
   VitalWireDelay (LEVEL0_ipd, LEVEL0, VitalExtendToFillDelay(tipd_LEVEL0));
   VitalWireDelay (LEVEL1_ipd, LEVEL1, VitalExtendToFillDelay(tipd_LEVEL1));
   VitalWireDelay (LEVEL2_ipd, LEVEL2, VitalExtendToFillDelay(tipd_LEVEL2));
   VitalWireDelay (LEVEL3_ipd, LEVEL3, VitalExtendToFillDelay(tipd_LEVEL3));
   VitalWireDelay (LEVEL4_ipd, LEVEL4, VitalExtendToFillDelay(tipd_LEVEL4));
   VitalWireDelay (LEVEL5_ipd, LEVEL5, VitalExtendToFillDelay(tipd_LEVEL5));
   VitalWireDelay (LEVEL6_ipd, LEVEL6, VitalExtendToFillDelay(tipd_LEVEL6));
   VitalWireDelay (LEVEL7_ipd, LEVEL7, VitalExtendToFillDelay(tipd_LEVEL7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RESET_ipd, RESET, VitalExtendToFillDelay(tipd_RESET));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

   ---------------------------------------------------------------
   --                  Behavior Section                         --
   ---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);

    VITALBehavior : process (
                          LEVEL0_ipd, LEVEL1_ipd, LEVEL2_ipd, LEVEL3_ipd, LEVEL4_ipd, LEVEL5_ipd, LEVEL6_ipd, LEVEL7_ipd, 
                          LGDEP0_ipd, LGDEP1_ipd, LGDEP2_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd, RESET_ipd
                          )

     -- some internal veriable declaration
     variable RAM_di_int   : std_logic_vector(8 downto 0);
     variable memory_array : MEM_TYPE  := (others =>(others => 'X'));
     variable do_par       : std_logic := 'X';
     variable tmp_par      : std_logic := 'X';
     variable tmp_par2     : std_logic := 'X';
     variable wpe_var      : std_logic := 'X';
     variable temp         : integer   := 0;
     variable thresh       : integer   := 0;
     variable depth        : integer   := 0;
     variable WADDR        : integer   := 0;
     variable WADDR_wrap   : integer   := 0;
     variable RADDR        : integer   := 0;
     variable RADDR_wrap   : integer   := 0;

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     --  Read Timing Check Results
     variable PeriodData_RESET           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET                : X01                 := '0';
     variable PeriodData_RDB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RDB                  : X01                 := '0';
     variable PeriodData_RBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RBLKB                : X01                 := '0';
     variable PeriodData_WRB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WRB                  : X01                 := '0';
     variable PeriodData_WBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WBLKB                : X01                 := '0';
     variable Tviol_DI0_WRB_posedge      : X01                 := '0';
     variable TmDt_DI0_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI0_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WRB_posedge      : X01                 := '0';
     variable TmDt_DI1_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI1_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WRB_posedge      : X01                 := '0';
     variable TmDt_DI2_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI2_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WRB_posedge      : X01                 := '0';
     variable TmDt_DI3_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI3_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WRB_posedge      : X01                 := '0';
     variable TmDt_DI4_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI4_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WRB_posedge      : X01                 := '0';
     variable TmDt_DI5_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI5_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WRB_posedge      : X01                 := '0';
     variable TmDt_DI6_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI6_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WRB_posedge      : X01                 := '0';
     variable TmDt_DI7_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI7_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WRB_posedge      : X01                 := '0';
     variable TmDt_DI8_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI8_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_RESET_posedge    : X01                 := '0';
     variable TmDt_WRB_RESET_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_RESET_posedge  : X01                 := '0';
     variable TmDt_WBLKB_RESET_posedge   : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results


     variable DO0_zd   : std_ulogic;
     variable DO1_zd   : std_ulogic;
     variable DO2_zd   : std_ulogic;
     variable DO3_zd   : std_ulogic;
     variable DO4_zd   : std_ulogic;
     variable DO5_zd   : std_ulogic;
     variable DO6_zd   : std_ulogic;
     variable DO7_zd   : std_ulogic;
     variable DO8_zd   : std_ulogic;
     variable RPE_zd   : std_ulogic;
     variable WPE_zd   : std_ulogic;
     variable DOS_zd   : std_ulogic;
     variable FULL_zd  : std_ulogic;
     variable EMPTY_zd : std_ulogic;
     variable EQTH_zd  : std_ulogic;
     variable GEQTH_zd : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData   : VitalGlitchDataType;
     variable DO1_GlitchData   : VitalGlitchDataType;
     variable DO2_GlitchData   : VitalGlitchDataType;
     variable DO3_GlitchData   : VitalGlitchDataType;
     variable DO4_GlitchData   : VitalGlitchDataType;
     variable DO5_GlitchData   : VitalGlitchDataType;
     variable DO6_GlitchData   : VitalGlitchDataType;
     variable DO7_GlitchData   : VitalGlitchDataType;
     variable DO8_GlitchData   : VitalGlitchDataType;
     variable RPE_GlitchData   : VitalGlitchDataType;
     variable WPE_GlitchData   : VitalGlitchDataType;
     variable DOS_GlitchData   : VitalGlitchDataType;
     variable FULL_GlitchData  : VitalGlitchDataType;
     variable EMPTY_GlitchData : VitalGlitchDataType;
     variable EQTH_GlitchData  : VitalGlitchDataType;
     variable GEQTH_GlitchData : VitalGlitchDataType;

     -- last value variables
     variable RBint_previous   : std_ulogic := 'X';
     variable WBint_previous   : std_ulogic := 'X';
     variable DIS_previous     : std_ulogic := 'X';
     variable RESET_previous   : std_ulogic := 'X';
     variable RESET_delayed    : std_ulogic := 'X';
     variable PARODD_previous  : std_ulogic := 'X';
     variable PARODD_delayed   : std_ulogic := 'X';
     variable DI0_delayed      : std_ulogic := 'X';
     variable DI1_delayed      : std_ulogic := 'X';
     variable DI2_delayed      : std_ulogic := 'X';
     variable DI3_delayed      : std_ulogic := 'X';
     variable DI4_delayed      : std_ulogic := 'X';
     variable DI5_delayed      : std_ulogic := 'X';
     variable DI6_delayed      : std_ulogic := 'X';
     variable DI7_delayed      : std_ulogic := 'X';
     variable DI8_delayed      : std_ulogic := 'X';
     variable DI0_previous     : std_ulogic := 'X';
     variable DI1_previous     : std_ulogic := 'X';
     variable DI2_previous     : std_ulogic := 'X';
     variable DI3_previous     : std_ulogic := 'X';
     variable DI4_previous     : std_ulogic := 'X';
     variable DI5_previous     : std_ulogic := 'X';
     variable DI6_previous     : std_ulogic := 'X';
     variable DI7_previous     : std_ulogic := 'X';
     variable DI8_previous     : std_ulogic := 'X';
     variable LGDEP0_delayed   : std_ulogic := 'X';
     variable LGDEP1_delayed   : std_ulogic := 'X';
     variable LGDEP2_delayed   : std_ulogic := 'X';
     variable LGDEP0_previous  : std_ulogic := 'X';
     variable LGDEP1_previous  : std_ulogic := 'X';
     variable LGDEP2_previous  : std_ulogic := 'X';
     variable LEVEL0_delayed   : std_ulogic := 'X';
     variable LEVEL1_delayed   : std_ulogic := 'X';
     variable LEVEL2_delayed   : std_ulogic := 'X';
     variable LEVEL3_delayed   : std_ulogic := 'X';
     variable LEVEL4_delayed   : std_ulogic := 'X';
     variable LEVEL5_delayed   : std_ulogic := 'X';
     variable LEVEL6_delayed   : std_ulogic := 'X';
     variable LEVEL7_delayed   : std_ulogic := 'X';
     variable LEVEL0_previous  : std_ulogic := 'X';
     variable LEVEL1_previous  : std_ulogic := 'X';
     variable LEVEL2_previous  : std_ulogic := 'X';
     variable LEVEL3_previous  : std_ulogic := 'X';
     variable LEVEL4_previous  : std_ulogic := 'X';
     variable LEVEL5_previous  : std_ulogic := 'X';
     variable LEVEL6_previous  : std_ulogic := 'X';
     variable LEVEL7_previous  : std_ulogic := 'X';

     variable WB_initialized   : Boolean := False; 
     -- True = WB_int falling edge occured.  
     -- Must occur before first write after RESET.
     
     -- Special variables to control flags
     variable hold_empty_low   : integer := 0;
     variable hold_eqth_high   : integer := 0;
     variable hold_geqth_high  : integer := 0;

 begin -- process VITALBehavior

 if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

      VitalPeriodPulseCheck ( Pviol_RDB,
                              PeriodData_RDB,
                              RDB_ipd, "RDB",
                              0.0 ns,
                              tperiod_RDB,
                              tpw_RDB_posedge,
                              tpw_RDB_negedge,
                              (TO_X01(RBLKB) = '0') AND (TO_X01(RESET ) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9AA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RBLKB,
                              PeriodData_RBLKB,
                              RBLKB_ipd, "RBLKB",
                              0.0 ns,
                              tperiod_RBLKB,
                              tpw_RBLKB_posedge,
                              tpw_RBLKB_negedge,
                              (TO_X01(RDB) = '0') AND (TO_X01(RESET ) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9AA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RESET,
                              PeriodData_RESET,
                              RESET_ipd, "RESET",
                              0.0 ns,
                              tpw_RESET_negedge,
                              0.0 ns,
                              tpw_RESET_negedge,
                              True,
                              InstancePath & "/FIFO256x9AA",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

   -- setup /hold check for WRB/WBLKB to RESET signal ;
       VitalSetupHoldCheck ( Tviol_WRB_RESET_posedge,
                             TmDt_WRB_RESET_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             tsetup_WRB_RESET_posedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             thold_WRB_RESET_negedge_posedge,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_RESET_posedge,
                             TmDt_WBLKB_RESET_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             tsetup_WBLKB_RESET_posedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             thold_WBLKB_RESET_negedge_posedge,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_posedge_posedge,
                             tsetup_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_posedge_posedge,
                             tsetup_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_posedge_posedge,
                             tsetup_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_posedge_posedge,
                             tsetup_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_posedge_posedge,
                             tsetup_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_posedge_posedge,
                             tsetup_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_posedge_posedge,
                             tsetup_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_posedge_posedge,
                             tsetup_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_posedge_posedge,
                             tsetup_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_posedge_posedge,
                             tsetup_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_posedge_posedge,
                             tsetup_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_posedge_posedge,
                             tsetup_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_posedge_posedge,
                             tsetup_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_posedge_posedge,
                             tsetup_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_posedge_posedge,
                             tsetup_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_posedge_posedge,
                             tsetup_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_posedge_posedge,
                             tsetup_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_posedge_posedge,
                             tsetup_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AA",
                             True,
                             True,
                             WARNING
                             );
      VitalPeriodPulseCheck ( Pviol_WRB,
                              PeriodData_WRB,
                              WRB_ipd, "WRB",
                              0.0 ns,
                              tperiod_WRB,
                              tpw_WRB_posedge,
                              tpw_WRB_negedge,
                              (TO_X01(WBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9AA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_WBLKB,
                              PeriodData_WBLKB,
                              WBLKB_ipd, "WBLKB",
                              0.0 ns,
                              tperiod_WBLKB,
                              tpw_WBLKB_posedge,
                              tpw_WBLKB_negedge,
                              (TO_X01(WRB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9AA",
                              True,
                              True,
                              WARNING
                              );
 end if;

   ------------------------------------------------------------
   --               FIFO RESET                               --
   ------------------------------------------------------------

   if ( RESET_ipd'event and RESET_ipd = '0' ) then
       WADDR           := 0;
       RADDR           := 0;
       WADDR_wrap      := 0;
       RADDR_wrap      := 0;
       FULL_zd         := '0';
       EMPTY_zd        := '1';
       EQTH_zd         := '0';
       GEQTH_zd        := '0';
       WPE_zd          := 'X';
       WB_initialized  := False;
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
   end if;

   if ( RESET_ipd'event and RESET_ipd = '1' ) then
     if ( TO_X01 ( WBint ) = '0' ) then
       EMPTY_zd        := '0';
       EQTH_zd         := '1';
       GEQTH_zd        := '1';
       hold_empty_low  := 1;
       hold_eqth_high  := 1;
       hold_geqth_high := 1;
     end if;
   end if;

   if ( WBint'event ) then
     hold_empty_low  := 0;
     hold_eqth_high  := 0;
     hold_geqth_high := 0;
   end if;

   ------------------------------------------------------------
   -- WPE output                                           -
   ------------------------------------------------------------

   if ( PARODD_ipd'EVENT ) then
     WPE_zd := not WPE_zd;
     RPE_zd := not RPE_zd;
   end if;

   ------------------------------------------------------------
   -- WPE generation block                            -
   ------------------------------------------------------------

     tmp_par := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;
     par_f <= tmp_par ;
     tmp_par2 := (tmp_par xor DI8_ipd);
     par_f2 <=  tmp_par2;

     if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
         ( TO_X01 ( DI8_ipd )    = 'X' ) or
         ( TO_X01 ( DI7_ipd )    = 'X' ) or
         ( TO_X01 ( DI6_ipd )    = 'X' ) or
         ( TO_X01 ( DI5_ipd )    = 'X' ) or
         ( TO_X01 ( DI4_ipd )    = 'X' ) or
         ( TO_X01 ( DI3_ipd )    = 'X' ) or
         ( TO_X01 ( DI2_ipd )    = 'X' ) or
         ( TO_X01 ( DI1_ipd )    = 'X' ) or
         ( TO_X01 ( DI0_ipd )    = 'X' )
        ) then
       wpe_var  :=  'X';
     else
       if ( tmp_par2 /= PARODD_ipd ) then
         wpe_var  :=  '1';
       else
         wpe_var  :=  '0';
       end if;
     end if;
     RAM_di_int(8) := DI8_ipd;
     WPE_zd := wpe_var;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

   if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
   end if; 

   -----------------------------------------------------------
   --    calculate the depth and levels                     --
   -----------------------------------------------------------

    temp :=((INT(LGDEP2_delayed)*4) + (INT(LGDEP1_delayed)*2) + 
           (INT(LGDEP0_delayed)*1));

    case temp is 
         when 0 => depth := 2;
         when 1 => depth := 4;
         when 2 => depth := 8;
         when 3 => depth := 16;
         when 4 => depth := 32;
         when 5 => depth := 64;
         when 6 => depth := 128;
         when 7 => depth := 256;
         when others => depth := 0;
    end case;
    
    -- threshold value

    thresh := (INT(LEVEL7_delayed)*128) + (INT(LEVEL6_delayed)*64) + 
               (INT(LEVEL5_delayed)*32) + (INT(LEVEL4_delayed)*16) + 
               (INT(LEVEL3_delayed)*8) + (INT(LEVEL2_delayed)*4) + 
               (INT(LEVEL1_delayed)*2) + (INT(LEVEL0_delayed)*1); 

    if ( thresh = 0 or thresh = 255 ) then
      assert false
        report " Illegal level configuration, LEVEL cannot be 0 or 255 "
        severity failure;
    end if;

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

    if ( WBint'event AND WBint = '0') then
      if ( TO_X01 ( RESET_ipd ) = '1' ) then
        WB_initialized := True;
      end if;
    end if;

    if ( WBint = '1' ) then
      null;
    elsif ( WBint = '0' ) AND ( TO_X01 ( RESET_ipd ) = '1' ) then
      if ( FULL_zd = '0' ) then 
        RAM_di_int ( 7 downto 0 ) := DI7_ipd & DI6_ipd & 
                                     DI5_ipd & DI4_ipd & 
                                     DI3_ipd & DI2_ipd & 
                                     DI1_ipd & DI0_ipd;
        memory_array(WADDR) := RAM_di_int;
      end if;
    else 
      null;
    end if;
    if (( WBint'event AND WBint = '1' ) AND 
        ( TO_X01 ( RESET_delayed ) = '1' ) AND
        ( WB_initialized )) then
      if ( FULL_zd = '0' ) then 
        if ( WADDR < depth - 1  ) then
          WADDR := WADDR + 1;
        elsif ( WADDR  = depth - 1 ) then
          WADDR := 0;
          WADDR_wrap := 1 - WADDR_wrap;
        end if;
        if ( WADDR = RADDR ) then
          if ( RADDR_wrap /= WADDR_wrap ) then
            FULL_zd := '1';
            EMPTY_zd :='0';
          end if;
        end if; 
        if ( WADDR /= RADDR ) then
          EMPTY_zd := '0';
        end if;
        if ( RADDR_wrap = WADDR_wrap ) then
          if ( WADDR - RADDR = thresh ) then
            EQTH_zd := '1';
          else 
            EQTH_zd := '0';
          end if;
          if ( WADDR - RADDR >= thresh ) then
            GEQTH_zd := '1';
          else 
            GEQTH_zd := '0';
          end if;
        else 
          if (( depth - RADDR + WADDR ) = thresh ) then
            EQTH_zd := '1';
          else 
            EQTH_zd := '0';
          end if;
          if ( depth - RADDR + WADDR >= thresh ) then
            GEQTH_zd := '1';
          else 
            GEQTH_zd := '0';
          end if;
        end if; 
      end if; -- FULL = 0
    end if; -- WBint went high


  --------------------------------------------------------------------
  --          FIFO READ SECTION........                             --
  --------------------------------------------------------------------

  if(TO_X01(RBint) = 'X') then 
    if(TO_X01(RESET_ipd) /= '0') then 
      if(TO_X01(RBint_previous) /= 'X') then
        assert false
        report ": RDB or RBLKB unknown"
        severity error;
      end if;
     end if;
  elsif ((RBint'event AND TO_X01(RBint) = '0') AND (TO_X01(RESET_ipd) /= '0')) then
     if(EMPTY_zd /= '1') then
           DO0_zd  := memory_array(RADDR)(0);
           DO1_zd  := memory_array(RADDR)(1);
           DO2_zd  := memory_array(RADDR)(2);
           DO3_zd  := memory_array(RADDR)(3);
           DO4_zd  := memory_array(RADDR)(4);
           DO5_zd  := memory_array(RADDR)(5);
           DO6_zd  := memory_array(RADDR)(6);
           DO7_zd  := memory_array(RADDR)(7);
           DO8_zd  := memory_array(RADDR)(8);
     if(RADDR <depth-1  ) then
        RADDR := RADDR + 1;
     else
        RADDR :=(RADDR +1) mod  depth;
        RADDR_wrap :=1 - RADDR_wrap;
     end if;
             do_par  :=DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR
                       DO3_zd XOR DO2_zd XOR DO1_zd XOR DO0_zd;
             par_f <= do_par;
             if (do_par = 'X') then
               RPE_zd := 'X';
             elsif (do_par /= PARODD_ipd) then
               RPE_zd := '1';
             else
               RPE_zd :=  '0';
             end if;
     end if;
  else 
   null;
  end if;
  if ((RBint'event and TO_X01(RBint) ='1') AND (TO_X01(RESET_ipd) /='0')) then
    if(RADDR = WADDR ) then
     if(RADDR_wrap = WADDR_wrap) then
       EMPTY_zd := '1';
       FULL_zd   :=  '0';
     end if;
    end if;
    if(RADDR /= WADDR ) then
     FULL_zd  := '0';
    end if;
     if(WADDR_wrap = RADDR_wrap ) then
      if((WADDR - RADDR) = thresh ) then
       EQTH_zd := '1';
      else
        EQTH_zd := '0';
      end if;
      if((WADDR - RADDR) >= thresh ) then
        GEQTH_zd := '1';
      else
        GEQTH_zd := '0';
      end if;
    else 
     if((depth + WADDR - RADDR) = thresh ) then
       EQTH_zd := '1';
     else
        EQTH_zd := '0';
     end if;
     if((depth + WADDR - RADDR) >= thresh ) then
       GEQTH_zd := '1';
     else
       GEQTH_zd := '0';
     end if;
    end if;
   end if;

   -- Mimic odd silicon flag behavior coming out of RESET with WB low
   
   if ( hold_empty_low = 1 ) then
     EMPTY_zd := '0';
   end if;

   if ( hold_eqth_high = 1 ) then
     EQTH_zd := '1';
   end if;

   -- If LEVEL greater than DEPTH then GEQTH mimics FULL
   
   if ( hold_geqth_high = 1 ) then
     GEQTH_zd := '1';
   else
     if ( thresh > depth ) then
       GEQTH_zd := FULL_zd;
     end if;
   end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       RBint_previous   := RBint;
       WBint_previous   := WBint;
       LGDEP0_previous  := LGDEP0_delayed;
       LGDEP0_delayed   := LGDEP0_ipd;
       LGDEP1_previous  := LGDEP1_delayed;
       LGDEP1_delayed   := LGDEP1_ipd;
       LGDEP2_previous  := LGDEP2_delayed;
       LGDEP2_delayed   := LGDEP2_ipd;
       LEVEL0_previous  := LEVEL0_delayed;
       LEVEL0_delayed   := LEVEL0_ipd;
       LEVEL1_previous  := LEVEL1_delayed;
       LEVEL1_delayed   := LEVEL1_ipd;
       LEVEL2_previous  := LEVEL2_delayed;
       LEVEL2_delayed   := LEVEL2_ipd;
       LEVEL3_previous  := LEVEL3_delayed;
       LEVEL3_delayed   := LEVEL3_ipd;
       LEVEL4_previous  := LEVEL4_delayed;
       LEVEL4_delayed   := LEVEL4_ipd;
       LEVEL5_previous  := LEVEL5_delayed;
       LEVEL5_delayed   := LEVEL5_ipd;
       LEVEL6_previous  := LEVEL6_delayed;
       LEVEL6_delayed   := LEVEL6_ipd;
       LEVEL7_previous  := LEVEL7_delayed;
       LEVEL7_delayed   := LEVEL7_ipd;
       PARODD_previous  := PARODD_delayed; 
       PARODD_delayed   := PARODD_ipd;
       RESET_previous   := RESET_delayed; 
       RESET_delayed    := RESET_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
             OutSignal     => DOS,
             GlitchData    => DOS_GlitchData,
             OutSignalName => "DOS",
             OutTemp       => DOS_zd,

             Paths =>   (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
           OutSignal     => WPE,
           GlitchData    => WPE_GlitchData,
           OutSignalName => "WPE",
           OutTemp       => WPE_zd,

           Paths =>   (0 => (DI0_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI0_WPE), true),
                       1 => (DI1_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI1_WPE), true),
                       2 => (DI2_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI2_WPE), true),
                       3 => (DI3_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI3_WPE), true),
                       4 => (DI4_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI4_WPE), true),
                       5 => (DI5_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI5_WPE), true),
                       6 => (DI6_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI6_WPE), true),
                       7 => (DI7_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI7_WPE), true),
                       8 => (DI8_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI8_WPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO0), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO0), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO1), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO1), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO2), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO2), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO3), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO3), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO4), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO4), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO5), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO5), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO6), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO6), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO7), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO7), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO8), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO8), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => RPE,
           GlitchData    => RPE_GlitchData,
           OutSignalName => "RPE",
           OutTemp       => RPE_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_RPE), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_RPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => FULL,
           GlitchData    => FULL_GlitchData,
           OutSignalName => "FULL",
           OutTemp       => FULL_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_FULL), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_FULL), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_FULL), true),
                       3 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_FULL), true),
                       4 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_FULL), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EMPTY,
           GlitchData    => EMPTY_GlitchData,
           OutSignalName => "EMPTY",
           OutTemp       => EMPTY_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EMPTY), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_EMPTY), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_EMPTY), true),
                       3 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_EMPTY), true),
                       4 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_EMPTY), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EQTH,
           GlitchData    => EQTH_GlitchData,
           OutSignalName => "EQTH",
           OutTemp       => EQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EQTH), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_EQTH), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_EQTH), true),
                       3 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_EQTH), true),
                       4 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_EQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => GEQTH,
           GlitchData    => GEQTH_GlitchData,
           OutSignalName => "GEQTH",
           OutTemp       => GEQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_GEQTH), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_GEQTH), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_GEQTH), true),
                       3 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_GEQTH), true),
                       4 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_GEQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );


   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

LIBRARY a500k;
USE a500k.all;

entity FIFO256x9AAP is 
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tpw_RDB_posedge         : VitalDelayType        := 0.000 ns;
 	tpw_RDB_negedge         : VitalDelayType        := 0.000 ns;
 	tperiod_RDB             : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_posedge       : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_negedge       : VitalDelayType        := 0.000 ns;
 	tperiod_RBLKB           : VitalDelayType        := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;

  	-- WB falling edge hold to RESETB   
 	thold_WRB_RESET_posedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_RESET_posedge_posedge             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_RESET_posedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RESET_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_WRB_RESET_negedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WBLKB_RESET_negedge_posedge             : VitalDelayType := 0.000 ns;
	tsetup_WRB_RESET_negedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_RESET_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                               : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                               : VitalDelayType := 0.000 ns;
 	tperiod_WRB                                   : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');


ATTRIBUTE VITAL_LEVEL0 OF FIFO256x9AAP : entity IS True ;
END FIFO256x9AAP;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of FIFO256x9AAP is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal LGDEP0_ipd : std_ulogic := 'X';
   signal LGDEP1_ipd : std_ulogic := 'X';
   signal LGDEP2_ipd : std_ulogic := 'X';
   signal LEVEL0_ipd : std_ulogic := 'X';
   signal LEVEL1_ipd : std_ulogic := 'X';
   signal LEVEL2_ipd : std_ulogic := 'X';
   signal LEVEL3_ipd : std_ulogic := 'X';
   signal LEVEL4_ipd : std_ulogic := 'X';
   signal LEVEL5_ipd : std_ulogic := 'X';
   signal LEVEL6_ipd : std_ulogic := 'X';
   signal LEVEL7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal RESET_ipd  : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

   -- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic := 'X';
   signal par_f2     : std_logic := 'X';

   signal WRITE_AT_PREV_EDGE : std_logic := '0';
   signal READ_AT_PREV_EDGE  : std_logic := '0';

   begin  --  VITAL_ACT

   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (LGDEP0_ipd, LGDEP0, VitalExtendToFillDelay(tipd_LGDEP0));
   VitalWireDelay (LGDEP1_ipd, LGDEP1, VitalExtendToFillDelay(tipd_LGDEP1));
   VitalWireDelay (LGDEP2_ipd, LGDEP2, VitalExtendToFillDelay(tipd_LGDEP2));
   VitalWireDelay (LEVEL0_ipd, LEVEL0, VitalExtendToFillDelay(tipd_LEVEL0));
   VitalWireDelay (LEVEL1_ipd, LEVEL1, VitalExtendToFillDelay(tipd_LEVEL1));
   VitalWireDelay (LEVEL2_ipd, LEVEL2, VitalExtendToFillDelay(tipd_LEVEL2));
   VitalWireDelay (LEVEL3_ipd, LEVEL3, VitalExtendToFillDelay(tipd_LEVEL3));
   VitalWireDelay (LEVEL4_ipd, LEVEL4, VitalExtendToFillDelay(tipd_LEVEL4));
   VitalWireDelay (LEVEL5_ipd, LEVEL5, VitalExtendToFillDelay(tipd_LEVEL5));
   VitalWireDelay (LEVEL6_ipd, LEVEL6, VitalExtendToFillDelay(tipd_LEVEL6));
   VitalWireDelay (LEVEL7_ipd, LEVEL7, VitalExtendToFillDelay(tipd_LEVEL7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RESET_ipd, RESET, VitalExtendToFillDelay(tipd_RESET));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

   ---------------------------------------------------------------
   --                  Behavior Section                         --
   ---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);

    VITALBehavior : process (
                          LEVEL0_ipd, LEVEL1_ipd, LEVEL2_ipd, LEVEL3_ipd, LEVEL4_ipd, LEVEL5_ipd, LEVEL6_ipd, LEVEL7_ipd, 
                          LGDEP0_ipd, LGDEP1_ipd, LGDEP2_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd, RESET_ipd
                          )

     -- some internal veriable declaration
     variable RAM_di_int   : std_logic_vector(8 downto 0);
     variable memory_array : MEM_TYPE  := (others =>(others => 'X'));
     variable do_par       : std_logic := 'X';
     variable tmp_par      : std_logic := 'X';
     variable tmp_par2     : std_logic := 'X';
     variable wpe_var      : std_logic := 'X';
     variable temp         : integer   := 0;
     variable thresh       : integer   := 0;
     variable depth        : integer   := 0;
     variable WADDR        : integer   := 0;
     variable WADDR_wrap   : integer   := 0;
     variable RADDR        : integer   := 0;
     variable RADDR_wrap   : integer   := 0;

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     --  Read Timing Check Results
     variable PeriodData_RESET           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET                : X01                 := '0';
     variable PeriodData_RDB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RDB                  : X01                 := '0';
     variable PeriodData_RBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RBLKB                : X01                 := '0';
     variable PeriodData_WRB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WRB                  : X01                 := '0';
     variable PeriodData_WBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WBLKB                : X01                 := '0';
     variable Tviol_DI0_WRB_posedge      : X01                 := '0';
     variable TmDt_DI0_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI0_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WRB_posedge      : X01                 := '0';
     variable TmDt_DI1_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI1_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WRB_posedge      : X01                 := '0';
     variable TmDt_DI2_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI2_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WRB_posedge      : X01                 := '0';
     variable TmDt_DI3_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI3_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WRB_posedge      : X01                 := '0';
     variable TmDt_DI4_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI4_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WRB_posedge      : X01                 := '0';
     variable TmDt_DI5_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI5_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WRB_posedge      : X01                 := '0';
     variable TmDt_DI6_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI6_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WRB_posedge      : X01                 := '0';
     variable TmDt_DI7_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI7_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WRB_posedge      : X01                 := '0';
     variable TmDt_DI8_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI8_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_RESET_posedge    : X01                 := '0';
     variable TmDt_WRB_RESET_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_RESET_posedge  : X01                 := '0';
     variable TmDt_WBLKB_RESET_posedge   : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results


     variable DO0_zd   : std_ulogic;
     variable DO1_zd   : std_ulogic;
     variable DO2_zd   : std_ulogic;
     variable DO3_zd   : std_ulogic;
     variable DO4_zd   : std_ulogic;
     variable DO5_zd   : std_ulogic;
     variable DO6_zd   : std_ulogic;
     variable DO7_zd   : std_ulogic;
     variable DO8_zd   : std_ulogic;
     variable RPE_zd   : std_ulogic;
     variable WPE_zd   : std_ulogic;
     variable DOS_zd   : std_ulogic;
     variable FULL_zd  : std_ulogic;
     variable EMPTY_zd : std_ulogic;
     variable EQTH_zd  : std_ulogic;
     variable GEQTH_zd : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData   : VitalGlitchDataType;
     variable DO1_GlitchData   : VitalGlitchDataType;
     variable DO2_GlitchData   : VitalGlitchDataType;
     variable DO3_GlitchData   : VitalGlitchDataType;
     variable DO4_GlitchData   : VitalGlitchDataType;
     variable DO5_GlitchData   : VitalGlitchDataType;
     variable DO6_GlitchData   : VitalGlitchDataType;
     variable DO7_GlitchData   : VitalGlitchDataType;
     variable DO8_GlitchData   : VitalGlitchDataType;
     variable DOS_GlitchData   : VitalGlitchDataType;
     variable FULL_GlitchData  : VitalGlitchDataType;
     variable EMPTY_GlitchData : VitalGlitchDataType;
     variable EQTH_GlitchData  : VitalGlitchDataType;
     variable GEQTH_GlitchData : VitalGlitchDataType;

     -- last value variables
     variable RBint_previous   : std_ulogic := 'X';
     variable WBint_previous   : std_ulogic := 'X';
     variable DIS_previous     : std_ulogic := 'X';
     variable RESET_previous   : std_ulogic := 'X';
     variable RESET_delayed    : std_ulogic := 'X';
     variable PARODD_previous  : std_ulogic := 'X';
     variable PARODD_delayed   : std_ulogic := 'X';
     variable DI0_delayed      : std_ulogic := 'X';
     variable DI1_delayed      : std_ulogic := 'X';
     variable DI2_delayed      : std_ulogic := 'X';
     variable DI3_delayed      : std_ulogic := 'X';
     variable DI4_delayed      : std_ulogic := 'X';
     variable DI5_delayed      : std_ulogic := 'X';
     variable DI6_delayed      : std_ulogic := 'X';
     variable DI7_delayed      : std_ulogic := 'X';
     variable DI8_delayed      : std_ulogic := 'X';
     variable DI0_previous     : std_ulogic := 'X';
     variable DI1_previous     : std_ulogic := 'X';
     variable DI2_previous     : std_ulogic := 'X';
     variable DI3_previous     : std_ulogic := 'X';
     variable DI4_previous     : std_ulogic := 'X';
     variable DI5_previous     : std_ulogic := 'X';
     variable DI6_previous     : std_ulogic := 'X';
     variable DI7_previous     : std_ulogic := 'X';
     variable DI8_previous     : std_ulogic := 'X';
     variable LGDEP0_delayed   : std_ulogic := 'X';
     variable LGDEP1_delayed   : std_ulogic := 'X';
     variable LGDEP2_delayed   : std_ulogic := 'X';
     variable LGDEP0_previous  : std_ulogic := 'X';
     variable LGDEP1_previous  : std_ulogic := 'X';
     variable LGDEP2_previous  : std_ulogic := 'X';
     variable LEVEL0_delayed   : std_ulogic := 'X';
     variable LEVEL1_delayed   : std_ulogic := 'X';
     variable LEVEL2_delayed   : std_ulogic := 'X';
     variable LEVEL3_delayed   : std_ulogic := 'X';
     variable LEVEL4_delayed   : std_ulogic := 'X';
     variable LEVEL5_delayed   : std_ulogic := 'X';
     variable LEVEL6_delayed   : std_ulogic := 'X';
     variable LEVEL7_delayed   : std_ulogic := 'X';
     variable LEVEL0_previous  : std_ulogic := 'X';
     variable LEVEL1_previous  : std_ulogic := 'X';
     variable LEVEL2_previous  : std_ulogic := 'X';
     variable LEVEL3_previous  : std_ulogic := 'X';
     variable LEVEL4_previous  : std_ulogic := 'X';
     variable LEVEL5_previous  : std_ulogic := 'X';
     variable LEVEL6_previous  : std_ulogic := 'X';
     variable LEVEL7_previous  : std_ulogic := 'X';

     variable WB_initialized   : Boolean := False; 
     -- True = WB_int falling edge occured.  
     -- Must occur before first write after RESET.

     -- Special variables to control flags
     variable hold_empty_low   : integer := 0;
     variable hold_eqth_high   : integer := 0;
     variable hold_geqth_high  : integer := 0;

 begin -- process VITALBehavior

 if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

      VitalPeriodPulseCheck ( Pviol_RDB,
                              PeriodData_RDB,
                              RDB_ipd, "RDB",
                              0.0 ns,
                              tperiod_RDB,
                              tpw_RDB_posedge,
                              tpw_RDB_negedge,
                              (TO_X01(RBLKB) = '0') AND (TO_X01(RESET ) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9AAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RBLKB,
                              PeriodData_RBLKB,
                              RBLKB_ipd, "RBLKB",
                              0.0 ns,
                              tperiod_RBLKB,
                              tpw_RBLKB_posedge,
                              tpw_RBLKB_negedge,
                              (TO_X01(RDB) = '0') AND (TO_X01(RESET ) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9AAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RESET,
                              PeriodData_RESET,
                              RESET_ipd, "RESET",
                              0.0 ns,
                              tpw_RESET_negedge,
                              0.0 ns,
                              tpw_RESET_negedge,
                              True,
                              InstancePath & "/FIFO256x9AAP",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

   -- setup /hold check for WRB/WBLKB to RESET signal ;
       VitalSetupHoldCheck ( Tviol_WRB_RESET_posedge,
                             TmDt_WRB_RESET_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             tsetup_WRB_RESET_posedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             thold_WRB_RESET_negedge_posedge,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_RESET_posedge,
                             TmDt_WBLKB_RESET_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             tsetup_WBLKB_RESET_posedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             thold_WBLKB_RESET_negedge_posedge,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_posedge_posedge,
                             tsetup_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_posedge_posedge,
                             tsetup_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_posedge_posedge,
                             tsetup_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_posedge_posedge,
                             tsetup_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_posedge_posedge,
                             tsetup_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_posedge_posedge,
                             tsetup_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_posedge_posedge,
                             tsetup_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_posedge_posedge,
                             tsetup_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_posedge_posedge,
                             tsetup_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_posedge_posedge,
                             tsetup_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_posedge_posedge,
                             tsetup_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_posedge_posedge,
                             tsetup_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_posedge_posedge,
                             tsetup_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_posedge_posedge,
                             tsetup_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_posedge_posedge,
                             tsetup_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_posedge_posedge,
                             tsetup_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_posedge_posedge,
                             tsetup_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_posedge_posedge,
                             tsetup_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AAP",
                             True,
                             True,
                             WARNING
                             );
      VitalPeriodPulseCheck ( Pviol_WRB,
                              PeriodData_WRB,
                              WRB_ipd, "WRB",
                              0.0 ns,
                              tperiod_WRB,
                              tpw_WRB_posedge,
                              tpw_WRB_negedge,
                              (TO_X01(WBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9AAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_WBLKB,
                              PeriodData_WBLKB,
                              WBLKB_ipd, "WBLKB",
                              0.0 ns,
                              tperiod_WBLKB,
                              tpw_WBLKB_posedge,
                              tpw_WBLKB_negedge,
                              (TO_X01(WRB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9AAP",
                              True,
                              True,
                              WARNING
                              );
 end if;

   ------------------------------------------------------------
   --               FIFO RESET                               --
   ------------------------------------------------------------

   if ( RESET_ipd'event and RESET_ipd = '0' ) then
       WADDR           := 0;
       RADDR           := 0;
       WADDR_wrap      := 0;
       RADDR_wrap      := 0;
       FULL_zd         := '0';
       EMPTY_zd        := '1';
       EQTH_zd         := '0';
       GEQTH_zd        := '0';
       WB_initialized  := False;
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
   end if;

   if ( RESET_ipd'event and RESET_ipd = '1' ) then
     if ( TO_X01 ( WBint ) = '0' ) then
       EMPTY_zd        := '0';
       EQTH_zd         := '1';
       GEQTH_zd        := '1';
       hold_empty_low  := 1;
       hold_eqth_high  := 1;
       hold_geqth_high := 1;
     end if;
   end if;

   if ( WBint'event ) then
     hold_empty_low  := 0;
     hold_eqth_high  := 0;
     hold_geqth_high := 0;
   end if;


   ------------------------------------------------------------
   --         WPE generating block                            -
   ------------------------------------------------------------

     tmp_par  := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;
     par_f  <= tmp_par ;
     if (tmp_par /= PARODD_ipd) then
        wpe_var  :=  '1';
     else
        wpe_var  :=  '0';
     end if;
     RAM_di_int(8) := wpe_var;
     WPE_zd := wpe_var;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

   if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
   end if; 

   -----------------------------------------------------------
   --    calculate the depth and levels                     --
   -----------------------------------------------------------

    temp :=((INT(LGDEP2_delayed)*4) + (INT(LGDEP1_delayed)*2) + 
           (INT(LGDEP0_delayed)*1));

    case temp is 
         when 0 => depth := 2;
         when 1 => depth := 4;
         when 2 => depth := 8;
         when 3 => depth := 16;
         when 4 => depth := 32;
         when 5 => depth := 64;
         when 6 => depth := 128;
         when 7 => depth := 256;
         when others => depth := 0;
    end case;

    -- thresh value

    thresh := (INT(LEVEL7_delayed)*128) + (INT(LEVEL6_delayed)*64) + 
               (INT(LEVEL5_delayed)*32) + (INT(LEVEL4_delayed)*16) + 
               (INT(LEVEL3_delayed)*8) + (INT(LEVEL2_delayed)*4) + 
               (INT(LEVEL1_delayed)*2) + (INT(LEVEL0_delayed)*1); 

    if ( thresh = 0 or thresh = 255 ) then
      assert false
        report " Illegal level configuration, LEVEL cannot be 0 or 255 "
        severity failure;
    end if;

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

    if ( WBint'event AND WBint = '0') then
      if ( TO_X01 ( RESET_ipd ) = '1' ) then
        WB_initialized := True;
      end if;
    end if;

    if(WBint = '1') then
        null;
    elsif(WBint = '0') AND (TO_X01(RESET_ipd) = '1') then
        if(FULL_zd = '0') then 
        RAM_di_int(7 downto 0) := DI7_ipd & DI6_ipd & 
                                   DI5_ipd & DI4_ipd & 
                                   DI3_ipd & DI2_ipd & 
                                   DI1_ipd & DI0_ipd;
         memory_array(WADDR) := RAM_di_int;
       end if;
    else 
      null;
    end if;
    if (( WBint'event AND WBint = '1' ) AND 
        ( TO_X01 ( RESET_delayed ) = '1' ) AND
        ( WB_initialized )) then
      if(FULL_zd = '0') then 
       if(WADDR <depth-1  ) then
           WADDR := WADDR + 1;
       elsif( WADDR  = depth-1) then
         WADDR := 0;
         WADDR_wrap := 1 - WADDR_wrap;
       end if;
       if(WADDR   = RADDR ) then
         if(RADDR_wrap /= WADDR_wrap) then
            FULL_zd := '1';
            EMPTY_zd :='0';
         end if;
       end if; 
         if(WADDR   /= RADDR ) then
          EMPTY_zd := '0';
         end if;
          if(RADDR_wrap = WADDR_wrap) then
            if(WADDR - RADDR = thresh ) then
               EQTH_zd := '1';
            else 
               EQTH_zd := '0';
            end if;
            if(WADDR - RADDR >= thresh ) then
                GEQTH_zd := '1';
            else 
                GEQTH_zd := '0';
            end if;
          else 
           if((depth -RADDR + WADDR) = thresh ) then
               EQTH_zd := '1';
           else 
               EQTH_zd := '0';
           end if;
           if(depth - RADDR + WADDR >= thresh ) then
                GEQTH_zd := '1';
           else 
                GEQTH_zd := '0';
           end if;
         end if; 
        end if;
      end if;


  --------------------------------------------------------------------
  --          FIFO READ SECTION........                             --
  --------------------------------------------------------------------

  if(TO_X01(RBint) = 'X') then 
    if(TO_X01(RESET_ipd) /= '0') then 
      if(TO_X01(RBint_previous) /= 'X') then
        assert false
        report ": RDB or RBLKB unknown"
        severity error;
      end if;
     end if;
  elsif ((RBint'event AND TO_X01(RBint) = '0') AND (TO_X01(RESET_ipd) /= '0')) then
     if(EMPTY_zd /= '1') then
           DO0_zd  := memory_array(RADDR)(0);
           DO1_zd  := memory_array(RADDR)(1);
           DO2_zd  := memory_array(RADDR)(2);
           DO3_zd  := memory_array(RADDR)(3);
           DO4_zd  := memory_array(RADDR)(4);
           DO5_zd  := memory_array(RADDR)(5);
           DO6_zd  := memory_array(RADDR)(6);
           DO7_zd  := memory_array(RADDR)(7);
           DO8_zd  := memory_array(RADDR)(8);
     if(RADDR <depth-1  ) then
        RADDR := RADDR + 1;
     else
        RADDR :=(RADDR +1) mod  depth;
        RADDR_wrap :=1 - RADDR_wrap;
     end if;
             do_par  :=DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR
                       DO3_zd XOR DO2_zd XOR DO1_zd XOR DO0_zd;
             par_f <= do_par;
             if (do_par = 'X') then
               RPE_zd := 'X';
             elsif (do_par /= PARODD_ipd) then
               RPE_zd := '1';
             else
               RPE_zd :=  '0';
             end if;
     end if;
  else 
   null;
  end if;
  if ((RBint'event and TO_X01(RBint) ='1') AND (TO_X01(RESET_ipd) /='0')) then
    if(RADDR = WADDR ) then
     if(RADDR_wrap = WADDR_wrap) then
       EMPTY_zd := '1';
       FULL_zd   :=  '0';
     end if;
    end if;
    if(RADDR /= WADDR ) then
     FULL_zd  := '0';
    end if;
     if(WADDR_wrap = RADDR_wrap ) then
      if((WADDR - RADDR) = thresh ) then
       EQTH_zd := '1';
      else
       EQTH_zd := '0';
      end if;
      if((WADDR - RADDR) >= thresh ) then
       GEQTH_zd := '1';
      else
       GEQTH_zd := '0';
      end if;
    else 
     if((depth + WADDR - RADDR) = thresh ) then
       EQTH_zd := '1';
     else
       EQTH_zd := '0';
     end if;
     if((depth + WADDR - RADDR) >= thresh ) then
       GEQTH_zd := '1';
     else
       GEQTH_zd := '0';
     end if;
    end if;
   end if;
   

   -- Mimic odd silicon flag behavior coming out of RESET with WB low
   
   if ( hold_empty_low = 1 ) then
     EMPTY_zd := '0';
   end if;

   if ( hold_eqth_high = 1 ) then
     EQTH_zd := '1';
   end if;

   -- If LEVEL greater than DEPTH then GEQTH mimics FULL
   
   if ( hold_geqth_high = 1 ) then
     GEQTH_zd := '1';
   else
     if ( thresh > depth ) then
       GEQTH_zd := FULL_zd;
     end if;
   end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       RBint_previous   := RBint;
       WBint_previous   := WBint;
       LGDEP0_previous  := LGDEP0_delayed;
       LGDEP0_delayed   := LGDEP0_ipd;
       LGDEP1_previous  := LGDEP1_delayed;
       LGDEP1_delayed   := LGDEP1_ipd;
       LGDEP2_previous  := LGDEP2_delayed;
       LGDEP2_delayed   := LGDEP2_ipd;
       LEVEL0_previous  := LEVEL0_delayed;
       LEVEL0_delayed   := LEVEL0_ipd;
       LEVEL1_previous  := LEVEL1_delayed;
       LEVEL1_delayed   := LEVEL1_ipd;
       LEVEL2_previous  := LEVEL2_delayed;
       LEVEL2_delayed   := LEVEL2_ipd;
       LEVEL3_previous  := LEVEL3_delayed;
       LEVEL3_delayed   := LEVEL3_ipd;
       LEVEL4_previous  := LEVEL4_delayed;
       LEVEL4_delayed   := LEVEL4_ipd;
       LEVEL5_previous  := LEVEL5_delayed;
       LEVEL5_delayed   := LEVEL5_ipd;
       LEVEL6_previous  := LEVEL6_delayed;
       LEVEL6_delayed   := LEVEL6_ipd;
       LEVEL7_previous  := LEVEL7_delayed;
       LEVEL7_delayed   := LEVEL7_ipd;
       PARODD_previous  := PARODD_delayed; 
       PARODD_delayed   := PARODD_ipd;
       RESET_previous   := RESET_delayed; 
       RESET_delayed    := RESET_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
             OutSignal     => DOS,
             GlitchData    => DOS_GlitchData,
             OutSignalName => "DOS",
             OutTemp       => DOS_zd,

             Paths =>   (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO0), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO0), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO1), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO1), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO2), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO2), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO3), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO3), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO4), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO4), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO5), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO5), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO6), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO6), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO7), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO7), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO8), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO8), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => FULL,
           GlitchData    => FULL_GlitchData,
           OutSignalName => "FULL",
           OutTemp       => FULL_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_FULL), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_FULL), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_FULL), true),
                       3 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_FULL), true),
                       4 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_FULL), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EMPTY,
           GlitchData    => EMPTY_GlitchData,
           OutSignalName => "EMPTY",
           OutTemp       => EMPTY_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EMPTY), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_EMPTY), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_EMPTY), true),
                       3 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_EMPTY), true),
                       4 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_EMPTY), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EQTH,
           GlitchData    => EQTH_GlitchData,
           OutSignalName => "EQTH",
           OutTemp       => EQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EQTH), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_EQTH), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_EQTH), true),
                       3 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_EQTH), true),
                       4 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_EQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => GEQTH,
           GlitchData    => GEQTH_GlitchData,
           OutSignalName => "GEQTH",
           OutTemp       => GEQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_GEQTH), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_GEQTH), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_GEQTH), true),
                       3 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_GEQTH), true),
                       4 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_GEQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );


   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

LIBRARY a500k;
USE a500k.all;
entity FIFO256x9ASR is 

   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI0_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI1_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI2_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI3_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI4_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI5_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI6_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI7_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI8_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;

  	-- WB falling edge hold to RESETB   
 	thold_WRB_RESET_posedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_RESET_posedge_posedge             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_RESET_posedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RESET_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_WRB_RESET_negedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WBLKB_RESET_negedge_posedge             : VitalDelayType := 0.000 ns;
	tsetup_WRB_RESET_negedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_RESET_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                               : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                               : VitalDelayType := 0.000 ns;
 	tperiod_WRB                                   : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        WPE    :  OUT STD_LOGIC := 'X';
        RPE    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');


ATTRIBUTE VITAL_LEVEL0 OF FIFO256x9ASR : entity IS True ;
END FIFO256x9ASR;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of FIFO256x9ASR is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal LGDEP0_ipd : std_ulogic := 'X';
   signal LGDEP1_ipd : std_ulogic := 'X';
   signal LGDEP2_ipd : std_ulogic := 'X';
   signal LEVEL0_ipd : std_ulogic := 'X';
   signal LEVEL1_ipd : std_ulogic := 'X';
   signal LEVEL2_ipd : std_ulogic := 'X';
   signal LEVEL3_ipd : std_ulogic := 'X';
   signal LEVEL4_ipd : std_ulogic := 'X';
   signal LEVEL5_ipd : std_ulogic := 'X';
   signal LEVEL6_ipd : std_ulogic := 'X';
   signal LEVEL7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal RESET_ipd  : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

   -- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic := 'X';
   signal par_f2     : std_logic := 'X';

   signal WRITE_AT_PREV_EDGE : std_logic := '0';
   signal READ_AT_PREV_EDGE  : std_logic := '0';

   begin  --  VITAL_ACT

   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (LGDEP0_ipd, LGDEP0, VitalExtendToFillDelay(tipd_LGDEP0));
   VitalWireDelay (LGDEP1_ipd, LGDEP1, VitalExtendToFillDelay(tipd_LGDEP1));
   VitalWireDelay (LGDEP2_ipd, LGDEP2, VitalExtendToFillDelay(tipd_LGDEP2));
   VitalWireDelay (LEVEL0_ipd, LEVEL0, VitalExtendToFillDelay(tipd_LEVEL0));
   VitalWireDelay (LEVEL1_ipd, LEVEL1, VitalExtendToFillDelay(tipd_LEVEL1));
   VitalWireDelay (LEVEL2_ipd, LEVEL2, VitalExtendToFillDelay(tipd_LEVEL2));
   VitalWireDelay (LEVEL3_ipd, LEVEL3, VitalExtendToFillDelay(tipd_LEVEL3));
   VitalWireDelay (LEVEL4_ipd, LEVEL4, VitalExtendToFillDelay(tipd_LEVEL4));
   VitalWireDelay (LEVEL5_ipd, LEVEL5, VitalExtendToFillDelay(tipd_LEVEL5));
   VitalWireDelay (LEVEL6_ipd, LEVEL6, VitalExtendToFillDelay(tipd_LEVEL6));
   VitalWireDelay (LEVEL7_ipd, LEVEL7, VitalExtendToFillDelay(tipd_LEVEL7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RESET_ipd, RESET, VitalExtendToFillDelay(tipd_RESET));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

   ---------------------------------------------------------------
   --                  Behavior Section                         --
   ---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);

    VITALBehavior : process (
                          LEVEL0_ipd, LEVEL1_ipd, LEVEL2_ipd, LEVEL3_ipd, LEVEL4_ipd, LEVEL5_ipd, LEVEL6_ipd, LEVEL7_ipd, 
                          LGDEP0_ipd, LGDEP1_ipd, LGDEP2_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd, RESET_ipd
                          )

     -- some internal veriable declaration
     variable RAM_di_int   : std_logic_vector(8 downto 0);
     variable memory_array : MEM_TYPE  := (others =>(others => 'X'));
     variable do_par       : std_logic := 'X';
     variable tmp_par      : std_logic := 'X';
     variable tmp_par2     : std_logic := 'X';
     variable wpe_var      : std_logic := 'X';
     variable temp         : integer   := 0;
     variable thresh       : integer   := 0;
     variable depth        : integer   := 0;
     variable WADDR        : integer   := 0;
     variable WADDR_wrap   : integer   := 0;
     variable RADDR        : integer   := 0;
     variable RADDR_wrap   : integer   := 0;

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     --  Read Timing Check Results
     variable PeriodData_RESET           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET                : X01                 := '0';
     variable Tviol_PARODD_RCLKS_posedge : X01                 := '0';
     variable TmDt_PARODD_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_RCLKS_posedge  : X01                 := '0';
     variable Tmkr_RESET_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable PeriodData_WRB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WRB                  : X01                 := '0';
     variable PeriodData_WBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WBLKB                : X01                 := '0';
     variable Tviol_DI0_WRB_posedge      : X01                 := '0';
     variable TmDt_DI0_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI0_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WRB_posedge      : X01                 := '0';
     variable TmDt_DI1_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI1_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WRB_posedge      : X01                 := '0';
     variable TmDt_DI2_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI2_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WRB_posedge      : X01                 := '0';
     variable TmDt_DI3_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI3_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WRB_posedge      : X01                 := '0';
     variable TmDt_DI4_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI4_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WRB_posedge      : X01                 := '0';
     variable TmDt_DI5_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI5_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WRB_posedge      : X01                 := '0';
     variable TmDt_DI6_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI6_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WRB_posedge      : X01                 := '0';
     variable TmDt_DI7_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI7_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WRB_posedge      : X01                 := '0';
     variable TmDt_DI8_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI8_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_RESET_posedge    : X01                 := '0';
     variable TmDt_WRB_RESET_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_RESET_posedge  : X01                 := '0';
     variable TmDt_WBLKB_RESET_posedge   : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results


     variable DO0_zd    : std_ulogic;
     variable DO1_zd    : std_ulogic;
     variable DO2_zd    : std_ulogic;
     variable DO3_zd    : std_ulogic;
     variable DO4_zd    : std_ulogic;
     variable DO5_zd    : std_ulogic;
     variable DO6_zd    : std_ulogic;
     variable DO7_zd    : std_ulogic;
     variable DO8_zd    : std_ulogic;
     variable RPE_zd    : std_ulogic;
     variable WPE_zd    : std_ulogic;
     variable DOS_zd    : std_ulogic;
     variable FULL_zd   : std_ulogic;
     variable EMPTY_zd  : std_ulogic;
     variable EQTH_zd   : std_ulogic;
     variable GEQTH_zd  : std_ulogic;
     variable EMPTY_tmp : std_ulogic;
     variable EQTH_tmp  : std_ulogic;
     variable GEQTH_tmp : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData   : VitalGlitchDataType;
     variable DO1_GlitchData   : VitalGlitchDataType;
     variable DO2_GlitchData   : VitalGlitchDataType;
     variable DO3_GlitchData   : VitalGlitchDataType;
     variable DO4_GlitchData   : VitalGlitchDataType;
     variable DO5_GlitchData   : VitalGlitchDataType;
     variable DO6_GlitchData   : VitalGlitchDataType;
     variable DO7_GlitchData   : VitalGlitchDataType;
     variable DO8_GlitchData   : VitalGlitchDataType;
     variable RPE_GlitchData   : VitalGlitchDataType;
     variable WPE_GlitchData   : VitalGlitchDataType;
     variable DOS_GlitchData   : VitalGlitchDataType;
     variable FULL_GlitchData  : VitalGlitchDataType;
     variable EMPTY_GlitchData : VitalGlitchDataType;
     variable EQTH_GlitchData  : VitalGlitchDataType;
     variable GEQTH_GlitchData : VitalGlitchDataType;

     -- last value variables
     variable RCLKS_previous   : std_ulogic := 'X';
     variable RBint_delayed    : std_ulogic := 'X';
     variable RBint_previous   : std_ulogic := 'X';
     variable WBint_previous   : std_ulogic := 'X';
     variable DIS_previous     : std_ulogic := 'X';
     variable RESET_previous   : std_ulogic := 'X';
     variable RESET_delayed    : std_ulogic := 'X';
     variable PARODD_previous  : std_ulogic := 'X';
     variable PARODD_delayed   : std_ulogic := 'X';
     variable DI0_delayed      : std_ulogic := 'X';
     variable DI1_delayed      : std_ulogic := 'X';
     variable DI2_delayed      : std_ulogic := 'X';
     variable DI3_delayed      : std_ulogic := 'X';
     variable DI4_delayed      : std_ulogic := 'X';
     variable DI5_delayed      : std_ulogic := 'X';
     variable DI6_delayed      : std_ulogic := 'X';
     variable DI7_delayed      : std_ulogic := 'X';
     variable DI8_delayed      : std_ulogic := 'X';
     variable DI0_previous     : std_ulogic := 'X';
     variable DI1_previous     : std_ulogic := 'X';
     variable DI2_previous     : std_ulogic := 'X';
     variable DI3_previous     : std_ulogic := 'X';
     variable DI4_previous     : std_ulogic := 'X';
     variable DI5_previous     : std_ulogic := 'X';
     variable DI6_previous     : std_ulogic := 'X';
     variable DI7_previous     : std_ulogic := 'X';
     variable DI8_previous     : std_ulogic := 'X';
     variable LGDEP0_delayed   : std_ulogic := 'X';
     variable LGDEP1_delayed   : std_ulogic := 'X';
     variable LGDEP2_delayed   : std_ulogic := 'X';
     variable LGDEP0_previous  : std_ulogic := 'X';
     variable LGDEP1_previous  : std_ulogic := 'X';
     variable LGDEP2_previous  : std_ulogic := 'X';
     variable LEVEL0_delayed   : std_ulogic := 'X';
     variable LEVEL1_delayed   : std_ulogic := 'X';
     variable LEVEL2_delayed   : std_ulogic := 'X';
     variable LEVEL3_delayed   : std_ulogic := 'X';
     variable LEVEL4_delayed   : std_ulogic := 'X';
     variable LEVEL5_delayed   : std_ulogic := 'X';
     variable LEVEL6_delayed   : std_ulogic := 'X';
     variable LEVEL7_delayed   : std_ulogic := 'X';
     variable LEVEL0_previous  : std_ulogic := 'X';
     variable LEVEL1_previous  : std_ulogic := 'X';
     variable LEVEL2_previous  : std_ulogic := 'X';
     variable LEVEL3_previous  : std_ulogic := 'X';
     variable LEVEL4_previous  : std_ulogic := 'X';
     variable LEVEL5_previous  : std_ulogic := 'X';
     variable LEVEL6_previous  : std_ulogic := 'X';
     variable LEVEL7_previous  : std_ulogic := 'X';

     --  Pipelined temporary results
     variable RPE_stg1         : std_ulogic := 'X';
     variable DO0_stg1         : std_ulogic := 'X';
     variable DO1_stg1         : std_ulogic := 'X';
     variable DO2_stg1         : std_ulogic := 'X';
     variable DO3_stg1         : std_ulogic := 'X';
     variable DO4_stg1         : std_ulogic := 'X';
     variable DO5_stg1         : std_ulogic := 'X';
     variable DO6_stg1         : std_ulogic := 'X';
     variable DO7_stg1         : std_ulogic := 'X';
     variable DO8_stg1         : std_ulogic := 'X';

     variable WB_initialized   : Boolean := False; 
     -- True = WB_int falling edge occured.  
     -- Must occur before first write after RESET.

     -- Special variables to control flags
     variable hold_empty_low   : integer := 0;
     variable hold_eqth_high   : integer := 0;
     variable hold_geqth_high  : integer := 0;

 begin -- process VITALBehavior

 if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

  -- recovery / removal check for RCLKS to RESET signal ;
       VitalRecoveryRemovalCheck ( Tviol_RESET_RCLKS_posedge,
                             Tmkr_RESET_RCLKS_posedge,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             trecovery_RESET_RCLKS_posedge_negedge,
                             thold_RESET_RCLKS_posedge_posedge,
                             TRUE,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'), 
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             TRUE,
                             TRUE,
                             WARNING
                             );

   -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             ((TO_X01(RBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             ((TO_X01(RDB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_PARODD_RCLKS_posedge,
                             TmDt_PARODD_RCLKS_posedge,
                             PARODD_ipd, "PARODD",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_PARODD_RCLKS_posedge_posedge,
                             tsetup_PARODD_RCLKS_negedge_posedge,
                             thold_PARODD_RCLKS_posedge_posedge,
                             thold_PARODD_RCLKS_negedge_posedge,
                             (TO_X01(RESET_ipd) = '1'),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (TO_X01(RDB) = '0') AND (TO_X01(RBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9ASR",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RESET,
                              PeriodData_RESET,
                              RESET_ipd, "RESET",
                              0.0 ns,
                              tpw_RESET_negedge,
                              0.0 ns,
                              tpw_RESET_negedge,
                              True,
                              InstancePath & "/FIFO256x9ASR",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

   -- setup /hold check for WRB/WBLKB to RESET signal ;
       VitalSetupHoldCheck ( Tviol_WRB_RESET_posedge,
                             TmDt_WRB_RESET_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             tsetup_WRB_RESET_posedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             thold_WRB_RESET_negedge_posedge,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_RESET_posedge,
                             TmDt_WBLKB_RESET_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             tsetup_WBLKB_RESET_posedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             thold_WBLKB_RESET_negedge_posedge,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_posedge_posedge,
                             tsetup_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_posedge_posedge,
                             tsetup_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_posedge_posedge,
                             tsetup_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_posedge_posedge,
                             tsetup_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_posedge_posedge,
                             tsetup_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_posedge_posedge,
                             tsetup_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_posedge_posedge,
                             tsetup_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_posedge_posedge,
                             tsetup_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_posedge_posedge,
                             tsetup_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_posedge_posedge,
                             tsetup_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_posedge_posedge,
                             tsetup_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_posedge_posedge,
                             tsetup_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_posedge_posedge,
                             tsetup_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_posedge_posedge,
                             tsetup_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_posedge_posedge,
                             tsetup_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_posedge_posedge,
                             tsetup_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_posedge_posedge,
                             tsetup_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_posedge_posedge,
                             tsetup_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASR",
                             True,
                             True,
                             WARNING
                             );
      VitalPeriodPulseCheck ( Pviol_WRB,
                              PeriodData_WRB,
                              WRB_ipd, "WRB",
                              0.0 ns,
                              tperiod_WRB,
                              tpw_WRB_posedge,
                              tpw_WRB_negedge,
                              (TO_X01(WBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9ASR",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_WBLKB,
                              PeriodData_WBLKB,
                              WBLKB_ipd, "WBLKB",
                              0.0 ns,
                              tperiod_WBLKB,
                              tpw_WBLKB_posedge,
                              tpw_WBLKB_negedge,
                              (TO_X01(WRB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9ASR",
                              True,
                              True,
                              WARNING
                              );
 end if;

   ------------------------------------------------------------
   --               FIFO RESET                               --
   ------------------------------------------------------------

   if(RESET_ipd'event AND RESET_ipd = '0') then
       WADDR      := 0;
       RADDR      := 0;
       WADDR_wrap := 0;
       RADDR_wrap := 0;
       FULL_zd    := '0';
       EMPTY_tmp  := '1';
       EQTH_tmp   := '0';
       GEQTH_tmp  := '0';
       READ_AT_PREV_EDGE <='0';
       WPE_zd     := 'X';
       WB_initialized := False;
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
   end if;

   if ( RESET_ipd'event and RESET_ipd = '1' ) then
     if ( TO_X01 ( WBint ) = '0' ) then
       EMPTY_zd        := '0';
       EQTH_zd         := '1';
       GEQTH_zd        := '1';
       hold_empty_low  := 1;
       hold_eqth_high  := 1;
       hold_geqth_high := 1;
     end if;
   end if;

   if ( WBint'event ) then
     hold_empty_low  := 0;
     hold_eqth_high  := 0;
     hold_geqth_high := 0;
   end if;

   ------------------------------------------------------------
   -- WPE output                                              -
   ------------------------------------------------------------

   if ( PARODD_ipd'EVENT ) then
     WPE_zd   := not WPE_zd;
     RPE_zd   := not RPE_zd;
     RPE_stg1 := not RPE_stg1;
   end if;

   ------------------------------------------------------------
   -- WPE generation block                                    -
   ------------------------------------------------------------

     tmp_par  := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;
     par_f  <= tmp_par ;
     tmp_par2 := (tmp_par xor DI8_ipd);
     par_f2  <=  tmp_par2;

     if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
         ( TO_X01 ( DI8_ipd )    = 'X' ) or
         ( TO_X01 ( DI7_ipd )    = 'X' ) or
         ( TO_X01 ( DI6_ipd )    = 'X' ) or
         ( TO_X01 ( DI5_ipd )    = 'X' ) or
         ( TO_X01 ( DI4_ipd )    = 'X' ) or
         ( TO_X01 ( DI3_ipd )    = 'X' ) or
         ( TO_X01 ( DI2_ipd )    = 'X' ) or
         ( TO_X01 ( DI1_ipd )    = 'X' ) or
         ( TO_X01 ( DI0_ipd )    = 'X' )
        ) then
       wpe_var  :=  'X';
     else
       if ( tmp_par2 /= PARODD_ipd ) then
         wpe_var  :=  '1';
       else
         wpe_var  :=  '0';
       end if;
     end if;
     RAM_di_int(8) := DI8_ipd;
     WPE_zd := wpe_var;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

   if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
   end if; 

   -----------------------------------------------------------
   --    calculate the depth and levels                     --
   -----------------------------------------------------------

    temp :=((INT(LGDEP2_delayed)*4) + (INT(LGDEP1_delayed)*2) + 
           (INT(LGDEP0_delayed)*1));

    case temp is 
         when 0 => depth := 2;
         when 1 => depth := 4;
         when 2 => depth := 8;
         when 3 => depth := 16;
         when 4 => depth := 32;
         when 5 => depth := 64;
         when 6 => depth := 128;
         when 7 => depth := 256;
         when others => depth := 0;
    end case;

    -- thresh value

    thresh := (INT(LEVEL7_delayed)*128) + (INT(LEVEL6_delayed)*64) + 
               (INT(LEVEL5_delayed)*32) + (INT(LEVEL4_delayed)*16) + 
               (INT(LEVEL3_delayed)*8) + (INT(LEVEL2_delayed)*4) + 
               (INT(LEVEL1_delayed)*2) + (INT(LEVEL0_delayed)*1); 

    if ( thresh = 0 or thresh = 255 ) then
      assert false
        report " Illegal level configuration, LEVEL cannot be 0 or 255 "
        severity failure;
    end if;

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

    if ( WBint'event AND WBint = '0') then
      if ( TO_X01 ( RESET_ipd ) = '1' ) then
        WB_initialized := True;
      end if;
    end if;

    if(WBint = '1') then
        null;
    elsif(WBint = '0') AND (TO_X01(RESET_ipd) = '1') then
        if(FULL_zd = '0') then 
        RAM_di_int(7 downto 0) := DI7_ipd & DI6_ipd & 
                                   DI5_ipd & DI4_ipd & 
                                   DI3_ipd & DI2_ipd & 
                                   DI1_ipd & DI0_ipd;
         memory_array(WADDR) := RAM_di_int;
       end if;
    else 
      null;
    end if;
    if (( WBint'event AND WBint = '1' ) AND 
        ( TO_X01 ( RESET_delayed ) = '1' ) AND
        ( WB_initialized )) then
      if(FULL_zd = '0') then 
       if(WADDR <depth-1  ) then
           WADDR := WADDR + 1;
       elsif( WADDR  = depth-1) then
         WADDR := 0;
         WADDR_wrap := 1 - WADDR_wrap;
       end if;
       if(WADDR   = RADDR ) then
         if(RADDR_wrap /= WADDR_wrap) then
            FULL_zd := '1';
            EMPTY_tmp :='0';
         end if;
       end if; 
         if(WADDR   /= RADDR ) then
          EMPTY_tmp := '0';
         end if;
          if(RADDR_wrap = WADDR_wrap) then
            if(WADDR - RADDR = thresh ) then
               EQTH_tmp := '1';
            else 
               EQTH_tmp := '0';
            end if;
            if(WADDR - RADDR >= thresh ) then
                GEQTH_tmp := '1';
            else 
                GEQTH_tmp := '0';
            end if;
          else 
           if((depth -RADDR + WADDR) = thresh ) then
               EQTH_tmp := '1';
           else 
               EQTH_tmp := '0';
           end if;
           if(depth - RADDR + WADDR >= thresh ) then
                GEQTH_tmp := '1';
           else 
                GEQTH_tmp := '0';
           end if;
         end if; 
        end if;
      end if;


  --------------------------------------------------------------------
  --          FIFO READ SECTION........                             --
  --------------------------------------------------------------------

  if (TO_X01(RCLKS_ipd)='X') then
    if(RESET_ipd /= '0') then
    if(TO_X01(RBint_delayed) /= '1') then
      if(TO_X01(RCLKS_previous) /= 'X') then
        assert false
        report ": RCLK unknown"
        severity Error;
        DO0_zd  := 'X';
        DO1_zd  := 'X';
        DO2_zd  := 'X';
        DO3_zd  := 'X';
        DO4_zd  := 'X';
        DO5_zd  := 'X';
        DO6_zd  := 'X';
        DO7_zd  := 'X';
        DO8_zd  := 'X';
      end if;
     end if;
    end if;
   elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='1') AND (TO_X01(RESET_delayed) = '1')) then
     DO0_zd := DO0_stg1;
     DO1_zd := DO1_stg1;
     DO2_zd := DO2_stg1;
     DO3_zd := DO3_stg1;
     DO4_zd := DO4_stg1;
     DO5_zd := DO5_stg1;
     DO6_zd := DO6_stg1;
     DO7_zd := DO7_stg1;
     DO8_zd := DO8_stg1;
     RPE_zd := RPE_stg1;
     READ_AT_PREV_EDGE <='0';
     case (TO_X01(RBint_delayed)) is
        when '1' =>
                null;
        when '0' =>
         if(TO_X01(EMPTY_zd) /= '1') then 
           DO0_stg1  := memory_array(RADDR)(0);
           DO1_stg1  := memory_array(RADDR)(1);
           DO2_stg1  := memory_array(RADDR)(2);
           DO3_stg1  := memory_array(RADDR)(3);
           DO4_stg1  := memory_array(RADDR)(4);
           DO5_stg1  := memory_array(RADDR)(5);
           DO6_stg1  := memory_array(RADDR)(6);
           DO7_stg1  := memory_array(RADDR)(7);
           DO8_stg1  := memory_array(RADDR)(8);
           READ_AT_PREV_EDGE <='1';
           if(RADDR <depth-1  ) then
             RADDR := RADDR + 1;
           else
             RADDR :=(RADDR +1) mod  depth;
             RADDR_wrap :=1 - RADDR_wrap;
           end if;
      do_par  := DO8_stg1 XOR DO7_stg1 XOR DO6_stg1 XOR DO5_stg1 XOR DO4_stg1 XOR DO3_stg1 XOR
                 DO2_stg1 XOR DO1_stg1 XOR DO0_stg1;
            par_f <= do_par;
            if (do_par = 'X') then
             RPE_stg1 := 'X';
            elsif (do_par /= PARODD_delayed) then
             RPE_stg1  :=  '1';
            else
             RPE_stg1  :=  '0';
            end if;
         end if;
     when others =>
       if (TO_X01(RBint_previous) /= 'X') then
        assert false
        report ": RDB or RBLKB unknown"
        severity Error;
        end if;
           DO0_stg1  := 'X';
           DO1_stg1  := 'X';
           DO2_stg1  := 'X';
           DO3_stg1  := 'X';
           DO4_stg1  := 'X';
           DO5_stg1  := 'X';
           DO6_stg1  := 'X';
           DO7_stg1  := 'X';
           DO8_stg1  := 'X';
     end case;
  elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='0') AND (TO_X01(RESET_delayed) = '1') AND (TO_X01(READ_AT_PREV_EDGE) = '1')) then
   READ_AT_PREV_EDGE <='0';
   if(RADDR = WADDR ) then
    if(RADDR_wrap = WADDR_wrap) then
       EMPTY_tmp := '1';
       FULL_zd  := '0';
    end if;
   end if;
   if(RADDR /= WADDR ) then
    FULL_zd  := '0';
   end if;
    if(WADDR_wrap = RADDR_wrap ) then
     if((WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((WADDR - RADDR) >= thresh  ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    else 
     if((depth + WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((depth + WADDR - RADDR) >= thresh ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    end if;
 else 
    null;
 end if;


   -- Mimic odd silicon flag behavior coming out of RESET with WB low
   
   if ( hold_empty_low = 1 ) then
     EMPTY_zd := '0';
   else
     EMPTY_zd := EMPTY_tmp;
   end if;

   if ( hold_eqth_high = 1 ) then
     EQTH_zd := '1';
   else
     EQTH_zd := EQTH_tmp;
   end if;

   -- If LEVEL greater than DEPTH then GEQTH mimics FULL
   
   if ( hold_geqth_high = 1 ) then
     GEQTH_zd := '1';
   else
     if ( thresh > depth ) then
       GEQTH_zd := FULL_zd;
     else
       GEQTH_zd := GEQTH_tmp;
     end if;
   end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       RCLKS_previous   := RCLKS_ipd;
       RBint_previous   := RBint_delayed;
       RBint_delayed    := RBint;
       WBint_previous   := WBint;
       LGDEP0_previous  := LGDEP0_delayed;
       LGDEP0_delayed   := LGDEP0_ipd;
       LGDEP1_previous  := LGDEP1_delayed;
       LGDEP1_delayed   := LGDEP1_ipd;
       LGDEP2_previous  := LGDEP2_delayed;
       LGDEP2_delayed   := LGDEP2_ipd;
       LEVEL0_previous  := LEVEL0_delayed;
       LEVEL0_delayed   := LEVEL0_ipd;
       LEVEL1_previous  := LEVEL1_delayed;
       LEVEL1_delayed   := LEVEL1_ipd;
       LEVEL2_previous  := LEVEL2_delayed;
       LEVEL2_delayed   := LEVEL2_ipd;
       LEVEL3_previous  := LEVEL3_delayed;
       LEVEL3_delayed   := LEVEL3_ipd;
       LEVEL4_previous  := LEVEL4_delayed;
       LEVEL4_delayed   := LEVEL4_ipd;
       LEVEL5_previous  := LEVEL5_delayed;
       LEVEL5_delayed   := LEVEL5_ipd;
       LEVEL6_previous  := LEVEL6_delayed;
       LEVEL6_delayed   := LEVEL6_ipd;
       LEVEL7_previous  := LEVEL7_delayed;
       LEVEL7_delayed   := LEVEL7_ipd;
       PARODD_previous  := PARODD_delayed; 
       PARODD_delayed   := PARODD_ipd;
       RESET_previous   := RESET_delayed; 
       RESET_delayed    := RESET_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
             OutSignal     => DOS,
             GlitchData    => DOS_GlitchData,
             OutSignalName => "DOS",
             OutTemp       => DOS_zd,

             Paths =>   (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
           OutSignal     => WPE,
           GlitchData    => WPE_GlitchData,
           OutSignalName => "WPE",
           OutTemp       => WPE_zd,

           Paths =>   (0 => (DI0_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI0_WPE), true),
                       1 => (DI1_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI1_WPE), true),
                       2 => (DI2_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI2_WPE), true),
                       3 => (DI3_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI3_WPE), true),
                       4 => (DI4_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI4_WPE), true),
                       5 => (DI5_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI5_WPE), true),
                       6 => (DI6_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI6_WPE), true),
                       7 => (DI7_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI7_WPE), true),
                       8 => (DI8_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI8_WPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO0), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO1), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO2), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO3), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO4), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO5), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO6), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO7), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO8), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => RPE,
           GlitchData    => RPE_GlitchData,
           OutSignalName => "RPE",
           OutTemp       => RPE_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_RPE), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_RPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => FULL,
           GlitchData    => FULL_GlitchData,
           OutSignalName => "FULL",
           OutTemp       => FULL_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_FULL), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_FULL), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_FULL), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_FULL), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EMPTY,
           GlitchData    => EMPTY_GlitchData,
           OutSignalName => "EMPTY",
           OutTemp       => EMPTY_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EMPTY), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_EMPTY), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_EMPTY), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EMPTY), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EQTH,
           GlitchData    => EQTH_GlitchData,
           OutSignalName => "EQTH",
           OutTemp       => EQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EQTH), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_EQTH), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_EQTH), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => GEQTH,
           GlitchData    => GEQTH_GlitchData,
           OutSignalName => "GEQTH",
           OutTemp       => GEQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_GEQTH), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_GEQTH), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_GEQTH), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_GEQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );


   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

LIBRARY a500k;
USE a500k.all;

entity FIFO256x9ASRP is 
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;

  	-- WB falling edge hold to RESETB   
 	thold_WRB_RESET_posedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_RESET_posedge_posedge             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_RESET_posedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RESET_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_WRB_RESET_negedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WBLKB_RESET_negedge_posedge             : VitalDelayType := 0.000 ns;
	tsetup_WRB_RESET_negedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_RESET_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                               : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                               : VitalDelayType := 0.000 ns;
 	tperiod_WRB                                   : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');


ATTRIBUTE VITAL_LEVEL0 OF FIFO256x9ASRP : entity IS True ;
END FIFO256x9ASRP;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of FIFO256x9ASRP is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal LGDEP0_ipd : std_ulogic := 'X';
   signal LGDEP1_ipd : std_ulogic := 'X';
   signal LGDEP2_ipd : std_ulogic := 'X';
   signal LEVEL0_ipd : std_ulogic := 'X';
   signal LEVEL1_ipd : std_ulogic := 'X';
   signal LEVEL2_ipd : std_ulogic := 'X';
   signal LEVEL3_ipd : std_ulogic := 'X';
   signal LEVEL4_ipd : std_ulogic := 'X';
   signal LEVEL5_ipd : std_ulogic := 'X';
   signal LEVEL6_ipd : std_ulogic := 'X';
   signal LEVEL7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal RESET_ipd  : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

   -- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic := 'X';
   signal par_f2     : std_logic := 'X';

   signal WRITE_AT_PREV_EDGE : std_logic := '0';
   signal READ_AT_PREV_EDGE  : std_logic := '0';

   begin  --  VITAL_ACT

   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (LGDEP0_ipd, LGDEP0, VitalExtendToFillDelay(tipd_LGDEP0));
   VitalWireDelay (LGDEP1_ipd, LGDEP1, VitalExtendToFillDelay(tipd_LGDEP1));
   VitalWireDelay (LGDEP2_ipd, LGDEP2, VitalExtendToFillDelay(tipd_LGDEP2));
   VitalWireDelay (LEVEL0_ipd, LEVEL0, VitalExtendToFillDelay(tipd_LEVEL0));
   VitalWireDelay (LEVEL1_ipd, LEVEL1, VitalExtendToFillDelay(tipd_LEVEL1));
   VitalWireDelay (LEVEL2_ipd, LEVEL2, VitalExtendToFillDelay(tipd_LEVEL2));
   VitalWireDelay (LEVEL3_ipd, LEVEL3, VitalExtendToFillDelay(tipd_LEVEL3));
   VitalWireDelay (LEVEL4_ipd, LEVEL4, VitalExtendToFillDelay(tipd_LEVEL4));
   VitalWireDelay (LEVEL5_ipd, LEVEL5, VitalExtendToFillDelay(tipd_LEVEL5));
   VitalWireDelay (LEVEL6_ipd, LEVEL6, VitalExtendToFillDelay(tipd_LEVEL6));
   VitalWireDelay (LEVEL7_ipd, LEVEL7, VitalExtendToFillDelay(tipd_LEVEL7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RESET_ipd, RESET, VitalExtendToFillDelay(tipd_RESET));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

   ---------------------------------------------------------------
   --                  Behavior Section                         --
   ---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);

    VITALBehavior : process (
                          LEVEL0_ipd, LEVEL1_ipd, LEVEL2_ipd, LEVEL3_ipd, LEVEL4_ipd, LEVEL5_ipd, LEVEL6_ipd, LEVEL7_ipd, 
                          LGDEP0_ipd, LGDEP1_ipd, LGDEP2_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd, RESET_ipd
                          )

     -- some internal veriable declaration
     variable RAM_di_int   : std_logic_vector(8 downto 0);
     variable memory_array : MEM_TYPE  := (others =>(others => 'X'));
     variable do_par       : std_logic := 'X';
     variable tmp_par      : std_logic := 'X';
     variable tmp_par2     : std_logic := 'X';
     variable wpe_var      : std_logic := 'X';
     variable temp         : integer   := 0;
     variable thresh       : integer   := 0;
     variable depth        : integer   := 0;
     variable WADDR        : integer   := 0;
     variable WADDR_wrap   : integer   := 0;
     variable RADDR        : integer   := 0;
     variable RADDR_wrap   : integer   := 0;

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     --  Read Timing Check Results
     variable PeriodData_RESET           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET                : X01                 := '0';
     variable Tviol_PARODD_RCLKS_posedge : X01                 := '0';
     variable TmDt_PARODD_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_RCLKS_posedge  : X01                 := '0';
     variable Tmkr_RESET_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable PeriodData_WRB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WRB                  : X01                 := '0';
     variable PeriodData_WBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WBLKB                : X01                 := '0';
     variable Tviol_DI0_WRB_posedge      : X01                 := '0';
     variable TmDt_DI0_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI0_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WRB_posedge      : X01                 := '0';
     variable TmDt_DI1_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI1_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WRB_posedge      : X01                 := '0';
     variable TmDt_DI2_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI2_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WRB_posedge      : X01                 := '0';
     variable TmDt_DI3_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI3_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WRB_posedge      : X01                 := '0';
     variable TmDt_DI4_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI4_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WRB_posedge      : X01                 := '0';
     variable TmDt_DI5_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI5_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WRB_posedge      : X01                 := '0';
     variable TmDt_DI6_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI6_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WRB_posedge      : X01                 := '0';
     variable TmDt_DI7_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI7_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WRB_posedge      : X01                 := '0';
     variable TmDt_DI8_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI8_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_RESET_posedge    : X01                 := '0';
     variable TmDt_WRB_RESET_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_RESET_posedge  : X01                 := '0';
     variable TmDt_WBLKB_RESET_posedge   : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results


     variable DO0_zd   : std_ulogic;
     variable DO1_zd   : std_ulogic;
     variable DO2_zd   : std_ulogic;
     variable DO3_zd   : std_ulogic;
     variable DO4_zd   : std_ulogic;
     variable DO5_zd   : std_ulogic;
     variable DO6_zd   : std_ulogic;
     variable DO7_zd   : std_ulogic;
     variable DO8_zd   : std_ulogic;
     variable RPE_zd   : std_ulogic;
     variable WPE_zd   : std_ulogic;
     variable DOS_zd   : std_ulogic;
     variable FULL_zd  : std_ulogic;
     variable EMPTY_zd : std_ulogic;
     variable EQTH_zd  : std_ulogic;
     variable GEQTH_zd : std_ulogic;
     variable EMPTY_tmp : std_ulogic;
     variable EQTH_tmp  : std_ulogic;
     variable GEQTH_tmp : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData   : VitalGlitchDataType;
     variable DO1_GlitchData   : VitalGlitchDataType;
     variable DO2_GlitchData   : VitalGlitchDataType;
     variable DO3_GlitchData   : VitalGlitchDataType;
     variable DO4_GlitchData   : VitalGlitchDataType;
     variable DO5_GlitchData   : VitalGlitchDataType;
     variable DO6_GlitchData   : VitalGlitchDataType;
     variable DO7_GlitchData   : VitalGlitchDataType;
     variable DO8_GlitchData   : VitalGlitchDataType;
     variable DOS_GlitchData   : VitalGlitchDataType;
     variable FULL_GlitchData  : VitalGlitchDataType;
     variable EMPTY_GlitchData : VitalGlitchDataType;
     variable EQTH_GlitchData  : VitalGlitchDataType;
     variable GEQTH_GlitchData : VitalGlitchDataType;

     -- last value variables
     variable RCLKS_previous   : std_ulogic := 'X';
     variable RBint_delayed    : std_ulogic := 'X';
     variable RBint_previous   : std_ulogic := 'X';
     variable WBint_previous   : std_ulogic := 'X';
     variable DIS_previous     : std_ulogic := 'X';
     variable RESET_previous   : std_ulogic := 'X';
     variable RESET_delayed    : std_ulogic := 'X';
     variable PARODD_previous  : std_ulogic := 'X';
     variable PARODD_delayed   : std_ulogic := 'X';
     variable DI0_delayed      : std_ulogic := 'X';
     variable DI1_delayed      : std_ulogic := 'X';
     variable DI2_delayed      : std_ulogic := 'X';
     variable DI3_delayed      : std_ulogic := 'X';
     variable DI4_delayed      : std_ulogic := 'X';
     variable DI5_delayed      : std_ulogic := 'X';
     variable DI6_delayed      : std_ulogic := 'X';
     variable DI7_delayed      : std_ulogic := 'X';
     variable DI8_delayed      : std_ulogic := 'X';
     variable DI0_previous     : std_ulogic := 'X';
     variable DI1_previous     : std_ulogic := 'X';
     variable DI2_previous     : std_ulogic := 'X';
     variable DI3_previous     : std_ulogic := 'X';
     variable DI4_previous     : std_ulogic := 'X';
     variable DI5_previous     : std_ulogic := 'X';
     variable DI6_previous     : std_ulogic := 'X';
     variable DI7_previous     : std_ulogic := 'X';
     variable DI8_previous     : std_ulogic := 'X';
     variable LGDEP0_delayed   : std_ulogic := 'X';
     variable LGDEP1_delayed   : std_ulogic := 'X';
     variable LGDEP2_delayed   : std_ulogic := 'X';
     variable LGDEP0_previous  : std_ulogic := 'X';
     variable LGDEP1_previous  : std_ulogic := 'X';
     variable LGDEP2_previous  : std_ulogic := 'X';
     variable LEVEL0_delayed   : std_ulogic := 'X';
     variable LEVEL1_delayed   : std_ulogic := 'X';
     variable LEVEL2_delayed   : std_ulogic := 'X';
     variable LEVEL3_delayed   : std_ulogic := 'X';
     variable LEVEL4_delayed   : std_ulogic := 'X';
     variable LEVEL5_delayed   : std_ulogic := 'X';
     variable LEVEL6_delayed   : std_ulogic := 'X';
     variable LEVEL7_delayed   : std_ulogic := 'X';
     variable LEVEL0_previous  : std_ulogic := 'X';
     variable LEVEL1_previous  : std_ulogic := 'X';
     variable LEVEL2_previous  : std_ulogic := 'X';
     variable LEVEL3_previous  : std_ulogic := 'X';
     variable LEVEL4_previous  : std_ulogic := 'X';
     variable LEVEL5_previous  : std_ulogic := 'X';
     variable LEVEL6_previous  : std_ulogic := 'X';
     variable LEVEL7_previous  : std_ulogic := 'X';

     --  Pipelined temporary results
     variable RPE_stg1         : std_ulogic := 'X';
     variable DO0_stg1         : std_ulogic := 'X';
     variable DO1_stg1         : std_ulogic := 'X';
     variable DO2_stg1         : std_ulogic := 'X';
     variable DO3_stg1         : std_ulogic := 'X';
     variable DO4_stg1         : std_ulogic := 'X';
     variable DO5_stg1         : std_ulogic := 'X';
     variable DO6_stg1         : std_ulogic := 'X';
     variable DO7_stg1         : std_ulogic := 'X';
     variable DO8_stg1         : std_ulogic := 'X';

     variable WB_initialized   : Boolean := False; 
     -- True = WB_int falling edge occured.  
     -- Must occur before first write after RESET.

     -- Special variables to control flags
     variable hold_empty_low   : integer := 0;
     variable hold_eqth_high   : integer := 0;
     variable hold_geqth_high  : integer := 0;

 begin -- process VITALBehavior

 if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

  -- recovery / removal check for RCLKS to RESET signal ;
       VitalRecoveryRemovalCheck ( Tviol_RESET_RCLKS_posedge,
                             Tmkr_RESET_RCLKS_posedge,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             trecovery_RESET_RCLKS_posedge_negedge,
                             thold_RESET_RCLKS_posedge_posedge,
                             TRUE,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'), 
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             TRUE,
                             TRUE,
                             WARNING
                             );

   -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             ((TO_X01(RBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             ((TO_X01(RDB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_PARODD_RCLKS_posedge,
                             TmDt_PARODD_RCLKS_posedge,
                             PARODD_ipd, "PARODD",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_PARODD_RCLKS_posedge_posedge,
                             tsetup_PARODD_RCLKS_negedge_posedge,
                             thold_PARODD_RCLKS_posedge_posedge,
                             thold_PARODD_RCLKS_negedge_posedge,
                             (TO_X01(RESET_ipd) = '1'),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (TO_X01(RDB) = '0') AND (TO_X01(RBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9ASRP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RESET,
                              PeriodData_RESET,
                              RESET_ipd, "RESET",
                              0.0 ns,
                              tpw_RESET_negedge,
                              0.0 ns,
                              tpw_RESET_negedge,
                              True,
                              InstancePath & "/FIFO256x9ASRP",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

   -- setup /hold check for WRB/WBLKB to RESET signal ;
       VitalSetupHoldCheck ( Tviol_WRB_RESET_posedge,
                             TmDt_WRB_RESET_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             tsetup_WRB_RESET_posedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             thold_WRB_RESET_negedge_posedge,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_RESET_posedge,
                             TmDt_WBLKB_RESET_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             tsetup_WBLKB_RESET_posedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             thold_WBLKB_RESET_negedge_posedge,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_posedge_posedge,
                             tsetup_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_posedge_posedge,
                             tsetup_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_posedge_posedge,
                             tsetup_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_posedge_posedge,
                             tsetup_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_posedge_posedge,
                             tsetup_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_posedge_posedge,
                             tsetup_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_posedge_posedge,
                             tsetup_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_posedge_posedge,
                             tsetup_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_posedge_posedge,
                             tsetup_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_posedge_posedge,
                             tsetup_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_posedge_posedge,
                             tsetup_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_posedge_posedge,
                             tsetup_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_posedge_posedge,
                             tsetup_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_posedge_posedge,
                             tsetup_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_posedge_posedge,
                             tsetup_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_posedge_posedge,
                             tsetup_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_posedge_posedge,
                             tsetup_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_posedge_posedge,
                             tsetup_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASRP",
                             True,
                             True,
                             WARNING
                             );
      VitalPeriodPulseCheck ( Pviol_WRB,
                              PeriodData_WRB,
                              WRB_ipd, "WRB",
                              0.0 ns,
                              tperiod_WRB,
                              tpw_WRB_posedge,
                              tpw_WRB_negedge,
                              (TO_X01(WBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9ASRP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_WBLKB,
                              PeriodData_WBLKB,
                              WBLKB_ipd, "WBLKB",
                              0.0 ns,
                              tperiod_WBLKB,
                              tpw_WBLKB_posedge,
                              tpw_WBLKB_negedge,
                              (TO_X01(WRB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9ASRP",
                              True,
                              True,
                              WARNING
                              );
 end if;

   ------------------------------------------------------------
   --               FIFO RESET                               --
   ------------------------------------------------------------

   if(RESET_ipd'event AND RESET_ipd = '0') then
       WADDR      := 0;
       RADDR      := 0;
       WADDR_wrap := 0;
       RADDR_wrap := 0;
       FULL_zd    := '0';
       EMPTY_tmp  := '1';
       EQTH_tmp   := '0';
       GEQTH_tmp  := '0';
       READ_AT_PREV_EDGE <='0';
       WB_initialized := False;
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
   end if;

   if ( RESET_ipd'event and RESET_ipd = '1' ) then
     if ( TO_X01 ( WBint ) = '0' ) then
       EMPTY_zd        := '0';
       EQTH_zd         := '1';
       GEQTH_zd        := '1';
       hold_empty_low  := 1;
       hold_eqth_high  := 1;
       hold_geqth_high := 1;
     end if;
   end if;

   if ( WBint'event ) then
     hold_empty_low  := 0;
     hold_eqth_high  := 0;
     hold_geqth_high := 0;
   end if;

   ------------------------------------------------------------
   --         WPE generating block                            -
   ------------------------------------------------------------

     tmp_par  := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;
     par_f  <= tmp_par ;
     if (tmp_par /= PARODD_ipd) then
        wpe_var  :=  '1';
     else
        wpe_var  :=  '0';
     end if;
     RAM_di_int(8) := wpe_var;
     WPE_zd := wpe_var;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

   if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
   end if; 

   -----------------------------------------------------------
   --    calculate the depth and levels                     --
   -----------------------------------------------------------

    temp :=((INT(LGDEP2_delayed)*4) + (INT(LGDEP1_delayed)*2) + 
           (INT(LGDEP0_delayed)*1));

    case temp is 
         when 0 => depth := 2;
         when 1 => depth := 4;
         when 2 => depth := 8;
         when 3 => depth := 16;
         when 4 => depth := 32;
         when 5 => depth := 64;
         when 6 => depth := 128;
         when 7 => depth := 256;
         when others => depth := 0;
    end case;

    -- thresh value

    thresh := (INT(LEVEL7_delayed)*128) + (INT(LEVEL6_delayed)*64) + 
               (INT(LEVEL5_delayed)*32) + (INT(LEVEL4_delayed)*16) + 
               (INT(LEVEL3_delayed)*8) + (INT(LEVEL2_delayed)*4) + 
               (INT(LEVEL1_delayed)*2) + (INT(LEVEL0_delayed)*1); 

    if ( thresh = 0 or thresh = 255 ) then
      assert false
        report " Illegal level configuration, LEVEL cannot be 0 or 255 "
        severity failure;
    end if;

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

    if ( WBint'event AND WBint = '0') then
      if ( TO_X01 ( RESET_ipd ) = '1' ) then
        WB_initialized := True;
      end if;
    end if;

    if(WBint = '1') then
        null;
    elsif(WBint = '0') AND (TO_X01(RESET_ipd) = '1') then
        if(FULL_zd = '0') then 
        RAM_di_int(7 downto 0) := DI7_ipd & DI6_ipd & 
                                   DI5_ipd & DI4_ipd & 
                                   DI3_ipd & DI2_ipd & 
                                   DI1_ipd & DI0_ipd;
         memory_array(WADDR) := RAM_di_int;
       end if;
    else 
      null;
    end if;
    if (( WBint'event AND WBint = '1' ) AND 
        ( TO_X01 ( RESET_delayed ) = '1' ) AND
        ( WB_initialized )) then
      if(FULL_zd = '0') then 
       if(WADDR <depth-1  ) then
           WADDR := WADDR + 1;
       elsif( WADDR  = depth-1) then
         WADDR := 0;
         WADDR_wrap := 1 - WADDR_wrap;
       end if;
       if(WADDR   = RADDR ) then
         if(RADDR_wrap /= WADDR_wrap) then
            FULL_zd := '1';
            EMPTY_tmp :='0';
         end if;
       end if; 
         if(WADDR   /= RADDR ) then
          EMPTY_tmp := '0';
         end if;
          if(RADDR_wrap = WADDR_wrap) then
            if(WADDR - RADDR = thresh ) then
               EQTH_tmp := '1';
            else 
               EQTH_tmp := '0';
            end if;
            if(WADDR - RADDR >= thresh ) then
                GEQTH_tmp := '1';
            else 
                GEQTH_tmp := '0';
            end if;
          else 
           if((depth -RADDR + WADDR) = thresh ) then
               EQTH_tmp := '1';
           else 
               EQTH_tmp := '0';
           end if;
           if(depth - RADDR + WADDR >= thresh ) then
                GEQTH_tmp := '1';
           else 
                GEQTH_tmp := '0';
           end if;
         end if; 
        end if;
      end if;


  --------------------------------------------------------------------
  --          FIFO READ SECTION........                             --
  --------------------------------------------------------------------

  if (TO_X01(RCLKS_ipd)='X') then
    if(RESET_ipd /= '0') then
    if(TO_X01(RBint_delayed) /= '1') then
      if(TO_X01(RCLKS_previous) /= 'X') then
        assert false
        report ": RCLK unknown"
        severity Error;
        DO0_zd  := 'X';
        DO1_zd  := 'X';
        DO2_zd  := 'X';
        DO3_zd  := 'X';
        DO4_zd  := 'X';
        DO5_zd  := 'X';
        DO6_zd  := 'X';
        DO7_zd  := 'X';
        DO8_zd  := 'X';
      end if;
     end if;
    end if;
   elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='1') AND (TO_X01(RESET_delayed) = '1')) then
     DO0_zd := DO0_stg1;
     DO1_zd := DO1_stg1;
     DO2_zd := DO2_stg1;
     DO3_zd := DO3_stg1;
     DO4_zd := DO4_stg1;
     DO5_zd := DO5_stg1;
     DO6_zd := DO6_stg1;
     DO7_zd := DO7_stg1;
     DO8_zd := DO8_stg1;
     RPE_zd := RPE_stg1;
     READ_AT_PREV_EDGE <='0';
     case (TO_X01(RBint_delayed)) is
        when '1' =>
                null;
        when '0' =>
         if(TO_X01(EMPTY_zd) /= '1') then 
           DO0_stg1  := memory_array(RADDR)(0);
           DO1_stg1  := memory_array(RADDR)(1);
           DO2_stg1  := memory_array(RADDR)(2);
           DO3_stg1  := memory_array(RADDR)(3);
           DO4_stg1  := memory_array(RADDR)(4);
           DO5_stg1  := memory_array(RADDR)(5);
           DO6_stg1  := memory_array(RADDR)(6);
           DO7_stg1  := memory_array(RADDR)(7);
           DO8_stg1  := memory_array(RADDR)(8);
           READ_AT_PREV_EDGE <='1';
           if(RADDR <depth-1  ) then
             RADDR := RADDR + 1;
           else
             RADDR :=(RADDR +1) mod  depth;
             RADDR_wrap :=1 - RADDR_wrap;
           end if;
      do_par  := DO8_stg1 XOR DO7_stg1 XOR DO6_stg1 XOR DO5_stg1 XOR DO4_stg1 XOR DO3_stg1 XOR
                 DO2_stg1 XOR DO1_stg1 XOR DO0_stg1;
            par_f <= do_par;
            if (do_par = 'X') then
             RPE_stg1 := 'X';
            elsif (do_par /= PARODD_delayed) then
             RPE_stg1  :=  '1';
            else
             RPE_stg1  :=  '0';
            end if;
         end if;
     when others =>
       if (TO_X01(RBint_previous) /= 'X') then
        assert false
        report ": RDB or RBLKB unknown"
        severity Error;
        end if;
           DO0_stg1  := 'X';
           DO1_stg1  := 'X';
           DO2_stg1  := 'X';
           DO3_stg1  := 'X';
           DO4_stg1  := 'X';
           DO5_stg1  := 'X';
           DO6_stg1  := 'X';
           DO7_stg1  := 'X';
           DO8_stg1  := 'X';
     end case;
  elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='0') AND (TO_X01(RESET_delayed) = '1') AND (TO_X01(READ_AT_PREV_EDGE) = '1')) then
   READ_AT_PREV_EDGE <='0';
   if(RADDR = WADDR ) then
    if(RADDR_wrap = WADDR_wrap) then
       EMPTY_tmp := '1';
       FULL_zd  := '0';
    end if;
   end if;
   if(RADDR /= WADDR ) then
    FULL_zd  := '0';
   end if;
    if(WADDR_wrap = RADDR_wrap ) then
     if((WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((WADDR - RADDR) >= thresh  ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    else 
     if((depth + WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((depth + WADDR - RADDR) >= thresh ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    end if;
 else 
    null;
 end if;


   -- Mimic odd silicon flag behavior coming out of RESET with WB low
   
   if ( hold_empty_low = 1 ) then
     EMPTY_zd := '0';
   else
     EMPTY_zd := EMPTY_tmp;
   end if;

   if ( hold_eqth_high = 1 ) then
     EQTH_zd := '1';
   else
     EQTH_zd := EQTH_tmp;
   end if;

   -- If LEVEL greater than DEPTH then GEQTH mimics FULL
   
   if ( hold_geqth_high = 1 ) then
     GEQTH_zd := '1';
   else
     if ( thresh > depth ) then
       GEQTH_zd := FULL_zd;
     else
       GEQTH_zd := GEQTH_tmp;
     end if;
   end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       RCLKS_previous   := RCLKS_ipd;
       RBint_previous   := RBint_delayed;
       RBint_delayed    := RBint;
       WBint_previous   := WBint;
       LGDEP0_previous  := LGDEP0_delayed;
       LGDEP0_delayed   := LGDEP0_ipd;
       LGDEP1_previous  := LGDEP1_delayed;
       LGDEP1_delayed   := LGDEP1_ipd;
       LGDEP2_previous  := LGDEP2_delayed;
       LGDEP2_delayed   := LGDEP2_ipd;
       LEVEL0_previous  := LEVEL0_delayed;
       LEVEL0_delayed   := LEVEL0_ipd;
       LEVEL1_previous  := LEVEL1_delayed;
       LEVEL1_delayed   := LEVEL1_ipd;
       LEVEL2_previous  := LEVEL2_delayed;
       LEVEL2_delayed   := LEVEL2_ipd;
       LEVEL3_previous  := LEVEL3_delayed;
       LEVEL3_delayed   := LEVEL3_ipd;
       LEVEL4_previous  := LEVEL4_delayed;
       LEVEL4_delayed   := LEVEL4_ipd;
       LEVEL5_previous  := LEVEL5_delayed;
       LEVEL5_delayed   := LEVEL5_ipd;
       LEVEL6_previous  := LEVEL6_delayed;
       LEVEL6_delayed   := LEVEL6_ipd;
       LEVEL7_previous  := LEVEL7_delayed;
       LEVEL7_delayed   := LEVEL7_ipd;
       PARODD_previous  := PARODD_delayed; 
       PARODD_delayed   := PARODD_ipd;
       RESET_previous   := RESET_delayed; 
       RESET_delayed    := RESET_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
             OutSignal     => DOS,
             GlitchData    => DOS_GlitchData,
             OutSignalName => "DOS",
             OutTemp       => DOS_zd,

             Paths =>   (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO0), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO1), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO2), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO3), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO4), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO5), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO6), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO7), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO8), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => FULL,
           GlitchData    => FULL_GlitchData,
           OutSignalName => "FULL",
           OutTemp       => FULL_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_FULL), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_FULL), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_FULL), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_FULL), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EMPTY,
           GlitchData    => EMPTY_GlitchData,
           OutSignalName => "EMPTY",
           OutTemp       => EMPTY_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EMPTY), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_EMPTY), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_EMPTY), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EMPTY), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EQTH,
           GlitchData    => EQTH_GlitchData,
           OutSignalName => "EQTH",
           OutTemp       => EQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EQTH), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_EQTH), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_EQTH), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => GEQTH,
           GlitchData    => GEQTH_GlitchData,
           OutSignalName => "GEQTH",
           OutTemp       => GEQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_GEQTH), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_GEQTH), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_GEQTH), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_GEQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );


   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

LIBRARY a500k;
USE a500k.all;

entity FIFO256x9AST is 
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI0_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI1_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI2_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI3_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI4_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI5_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI6_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI7_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_DI8_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;

  	-- WB falling edge hold to RESETB   
 	thold_WRB_RESET_posedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_RESET_posedge_posedge             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_RESET_posedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RESET_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_WRB_RESET_negedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WBLKB_RESET_negedge_posedge             : VitalDelayType := 0.000 ns;
	tsetup_WRB_RESET_negedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_RESET_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                               : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                               : VitalDelayType := 0.000 ns;
 	tperiod_WRB                                   : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        WPE    :  OUT STD_LOGIC := 'X';
        RPE    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');


ATTRIBUTE VITAL_LEVEL0 OF FIFO256x9AST : entity IS True ;
END FIFO256x9AST;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of FIFO256x9AST is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal LGDEP0_ipd : std_ulogic := 'X';
   signal LGDEP1_ipd : std_ulogic := 'X';
   signal LGDEP2_ipd : std_ulogic := 'X';
   signal LEVEL0_ipd : std_ulogic := 'X';
   signal LEVEL1_ipd : std_ulogic := 'X';
   signal LEVEL2_ipd : std_ulogic := 'X';
   signal LEVEL3_ipd : std_ulogic := 'X';
   signal LEVEL4_ipd : std_ulogic := 'X';
   signal LEVEL5_ipd : std_ulogic := 'X';
   signal LEVEL6_ipd : std_ulogic := 'X';
   signal LEVEL7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal RESET_ipd  : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

   -- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic := 'X';
   signal par_f2     : std_logic := 'X';

   signal WRITE_AT_PREV_EDGE : std_logic := '0';
   signal READ_AT_PREV_EDGE  : std_logic := '0';

   begin  --  VITAL_ACT

   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (LGDEP0_ipd, LGDEP0, VitalExtendToFillDelay(tipd_LGDEP0));
   VitalWireDelay (LGDEP1_ipd, LGDEP1, VitalExtendToFillDelay(tipd_LGDEP1));
   VitalWireDelay (LGDEP2_ipd, LGDEP2, VitalExtendToFillDelay(tipd_LGDEP2));
   VitalWireDelay (LEVEL0_ipd, LEVEL0, VitalExtendToFillDelay(tipd_LEVEL0));
   VitalWireDelay (LEVEL1_ipd, LEVEL1, VitalExtendToFillDelay(tipd_LEVEL1));
   VitalWireDelay (LEVEL2_ipd, LEVEL2, VitalExtendToFillDelay(tipd_LEVEL2));
   VitalWireDelay (LEVEL3_ipd, LEVEL3, VitalExtendToFillDelay(tipd_LEVEL3));
   VitalWireDelay (LEVEL4_ipd, LEVEL4, VitalExtendToFillDelay(tipd_LEVEL4));
   VitalWireDelay (LEVEL5_ipd, LEVEL5, VitalExtendToFillDelay(tipd_LEVEL5));
   VitalWireDelay (LEVEL6_ipd, LEVEL6, VitalExtendToFillDelay(tipd_LEVEL6));
   VitalWireDelay (LEVEL7_ipd, LEVEL7, VitalExtendToFillDelay(tipd_LEVEL7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RESET_ipd, RESET, VitalExtendToFillDelay(tipd_RESET));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

   ---------------------------------------------------------------
   --                  Behavior Section                         --
   ---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);

    VITALBehavior : process (
                          LEVEL0_ipd, LEVEL1_ipd, LEVEL2_ipd, LEVEL3_ipd, LEVEL4_ipd, LEVEL5_ipd, LEVEL6_ipd, LEVEL7_ipd, 
                          LGDEP0_ipd, LGDEP1_ipd, LGDEP2_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd, RESET_ipd
                          )

     -- some internal veriable declaration
     variable RAM_di_int   : std_logic_vector(8 downto 0);
     variable memory_array : MEM_TYPE  := (others =>(others => 'X'));
     variable do_par       : std_logic := 'X';
     variable tmp_par      : std_logic := 'X';
     variable tmp_par2     : std_logic := 'X';
     variable wpe_var      : std_logic := 'X';
     variable temp         : integer   := 0;
     variable thresh       : integer   := 0;
     variable depth        : integer   := 0;
     variable WADDR        : integer   := 0;
     variable WADDR_wrap   : integer   := 0;
     variable RADDR        : integer   := 0;
     variable RADDR_wrap   : integer   := 0;

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     --  Read Timing Check Results
     variable PeriodData_RESET           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET                : X01                 := '0';
     variable Tviol_PARODD_RCLKS_posedge : X01                 := '0';
     variable TmDt_PARODD_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_RCLKS_posedge  : X01                 := '0';
     variable Tmkr_RESET_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable PeriodData_WRB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WRB                  : X01                 := '0';
     variable PeriodData_WBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WBLKB                : X01                 := '0';
     variable Tviol_DI0_WRB_posedge      : X01                 := '0';
     variable TmDt_DI0_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI0_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WRB_posedge      : X01                 := '0';
     variable TmDt_DI1_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI1_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WRB_posedge      : X01                 := '0';
     variable TmDt_DI2_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI2_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WRB_posedge      : X01                 := '0';
     variable TmDt_DI3_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI3_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WRB_posedge      : X01                 := '0';
     variable TmDt_DI4_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI4_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WRB_posedge      : X01                 := '0';
     variable TmDt_DI5_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI5_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WRB_posedge      : X01                 := '0';
     variable TmDt_DI6_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI6_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WRB_posedge      : X01                 := '0';
     variable TmDt_DI7_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI7_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WRB_posedge      : X01                 := '0';
     variable TmDt_DI8_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI8_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_RESET_posedge    : X01                 := '0';
     variable TmDt_WRB_RESET_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_RESET_posedge  : X01                 := '0';
     variable TmDt_WBLKB_RESET_posedge   : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results


     variable DO0_zd   : std_ulogic;
     variable DO1_zd   : std_ulogic;
     variable DO2_zd   : std_ulogic;
     variable DO3_zd   : std_ulogic;
     variable DO4_zd   : std_ulogic;
     variable DO5_zd   : std_ulogic;
     variable DO6_zd   : std_ulogic;
     variable DO7_zd   : std_ulogic;
     variable DO8_zd   : std_ulogic;
     variable RPE_zd   : std_ulogic;
     variable WPE_zd   : std_ulogic;
     variable DOS_zd   : std_ulogic;
     variable FULL_zd  : std_ulogic;
     variable EMPTY_zd : std_ulogic;
     variable EQTH_zd  : std_ulogic;
     variable GEQTH_zd : std_ulogic;
     variable EMPTY_tmp : std_ulogic;
     variable EQTH_tmp  : std_ulogic;
     variable GEQTH_tmp : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData   : VitalGlitchDataType;
     variable DO1_GlitchData   : VitalGlitchDataType;
     variable DO2_GlitchData   : VitalGlitchDataType;
     variable DO3_GlitchData   : VitalGlitchDataType;
     variable DO4_GlitchData   : VitalGlitchDataType;
     variable DO5_GlitchData   : VitalGlitchDataType;
     variable DO6_GlitchData   : VitalGlitchDataType;
     variable DO7_GlitchData   : VitalGlitchDataType;
     variable DO8_GlitchData   : VitalGlitchDataType;
     variable RPE_GlitchData   : VitalGlitchDataType;
     variable WPE_GlitchData   : VitalGlitchDataType;
     variable DOS_GlitchData   : VitalGlitchDataType;
     variable FULL_GlitchData  : VitalGlitchDataType;
     variable EMPTY_GlitchData : VitalGlitchDataType;
     variable EQTH_GlitchData  : VitalGlitchDataType;
     variable GEQTH_GlitchData : VitalGlitchDataType;

     -- last value variables
     variable RCLKS_previous   : std_ulogic := 'X';
     variable RBint_delayed    : std_ulogic := 'X';
     variable RBint_previous   : std_ulogic := 'X';
     variable WBint_previous   : std_ulogic := 'X';
     variable DIS_previous     : std_ulogic := 'X';
     variable RESET_previous   : std_ulogic := 'X';
     variable RESET_delayed    : std_ulogic := 'X';
     variable PARODD_previous  : std_ulogic := 'X';
     variable PARODD_delayed   : std_ulogic := 'X';
     variable DI0_delayed      : std_ulogic := 'X';
     variable DI1_delayed      : std_ulogic := 'X';
     variable DI2_delayed      : std_ulogic := 'X';
     variable DI3_delayed      : std_ulogic := 'X';
     variable DI4_delayed      : std_ulogic := 'X';
     variable DI5_delayed      : std_ulogic := 'X';
     variable DI6_delayed      : std_ulogic := 'X';
     variable DI7_delayed      : std_ulogic := 'X';
     variable DI8_delayed      : std_ulogic := 'X';
     variable DI0_previous     : std_ulogic := 'X';
     variable DI1_previous     : std_ulogic := 'X';
     variable DI2_previous     : std_ulogic := 'X';
     variable DI3_previous     : std_ulogic := 'X';
     variable DI4_previous     : std_ulogic := 'X';
     variable DI5_previous     : std_ulogic := 'X';
     variable DI6_previous     : std_ulogic := 'X';
     variable DI7_previous     : std_ulogic := 'X';
     variable DI8_previous     : std_ulogic := 'X';
     variable LGDEP0_delayed   : std_ulogic := 'X';
     variable LGDEP1_delayed   : std_ulogic := 'X';
     variable LGDEP2_delayed   : std_ulogic := 'X';
     variable LGDEP0_previous  : std_ulogic := 'X';
     variable LGDEP1_previous  : std_ulogic := 'X';
     variable LGDEP2_previous  : std_ulogic := 'X';
     variable LEVEL0_delayed   : std_ulogic := 'X';
     variable LEVEL1_delayed   : std_ulogic := 'X';
     variable LEVEL2_delayed   : std_ulogic := 'X';
     variable LEVEL3_delayed   : std_ulogic := 'X';
     variable LEVEL4_delayed   : std_ulogic := 'X';
     variable LEVEL5_delayed   : std_ulogic := 'X';
     variable LEVEL6_delayed   : std_ulogic := 'X';
     variable LEVEL7_delayed   : std_ulogic := 'X';
     variable LEVEL0_previous  : std_ulogic := 'X';
     variable LEVEL1_previous  : std_ulogic := 'X';
     variable LEVEL2_previous  : std_ulogic := 'X';
     variable LEVEL3_previous  : std_ulogic := 'X';
     variable LEVEL4_previous  : std_ulogic := 'X';
     variable LEVEL5_previous  : std_ulogic := 'X';
     variable LEVEL6_previous  : std_ulogic := 'X';
     variable LEVEL7_previous  : std_ulogic := 'X';

     variable WB_initialized   : Boolean := False; 
     -- True = WB_int falling edge occured.  
     -- Must occur before first write after RESET.

     -- Special variables to control flags
     variable hold_empty_low   : integer := 0;
     variable hold_eqth_high   : integer := 0;
     variable hold_geqth_high  : integer := 0;

 begin -- process VITALBehavior

 if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

   -- recovery / removal check for RCLKS to RESET signal ;
       VitalRecoveryRemovalCheck ( Tviol_RESET_RCLKS_posedge,
                             Tmkr_RESET_RCLKS_posedge,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             trecovery_RESET_RCLKS_posedge_negedge,
                             thold_RESET_RCLKS_posedge_posedge,
                             TRUE,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'), 
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             TRUE,
                             TRUE,
                             WARNING
                             );

   -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             ((TO_X01(RBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             ((TO_X01(RDB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_PARODD_RCLKS_posedge,
                             TmDt_PARODD_RCLKS_posedge,
                             PARODD_ipd, "PARODD",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_PARODD_RCLKS_posedge_posedge,
                             tsetup_PARODD_RCLKS_negedge_posedge,
                             thold_PARODD_RCLKS_posedge_posedge,
                             thold_PARODD_RCLKS_negedge_posedge,
                             (TO_X01(RESET_ipd) = '1'),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (TO_X01(RDB) = '0') AND (TO_X01(RBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9AST",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RESET,
                              PeriodData_RESET,
                              RESET_ipd, "RESET",
                              0.0 ns,
                              tpw_RESET_negedge,
                              0.0 ns,
                              tpw_RESET_negedge,
                              True,
                              InstancePath & "/FIFO256x9AST",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

   -- setup /hold check for WRB/WBLKB to RESET signal ;
       VitalSetupHoldCheck ( Tviol_WRB_RESET_posedge,
                             TmDt_WRB_RESET_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             tsetup_WRB_RESET_posedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             thold_WRB_RESET_negedge_posedge,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_RESET_posedge,
                             TmDt_WBLKB_RESET_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             tsetup_WBLKB_RESET_posedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             thold_WBLKB_RESET_negedge_posedge,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_posedge_posedge,
                             tsetup_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_posedge_posedge,
                             tsetup_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_posedge_posedge,
                             tsetup_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_posedge_posedge,
                             tsetup_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_posedge_posedge,
                             tsetup_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_posedge_posedge,
                             tsetup_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_posedge_posedge,
                             tsetup_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_posedge_posedge,
                             tsetup_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_posedge_posedge,
                             tsetup_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_posedge_posedge,
                             tsetup_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_posedge_posedge,
                             tsetup_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_posedge_posedge,
                             tsetup_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_posedge_posedge,
                             tsetup_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_posedge_posedge,
                             tsetup_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_posedge_posedge,
                             tsetup_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_posedge_posedge,
                             tsetup_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_posedge_posedge,
                             tsetup_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_posedge_posedge,
                             tsetup_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9AST",
                             True,
                             True,
                             WARNING
                             );
      VitalPeriodPulseCheck ( Pviol_WRB,
                              PeriodData_WRB,
                              WRB_ipd, "WRB",
                              0.0 ns,
                              tperiod_WRB,
                              tpw_WRB_posedge,
                              tpw_WRB_negedge,
                              (TO_X01(WBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9AST",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_WBLKB,
                              PeriodData_WBLKB,
                              WBLKB_ipd, "WBLKB",
                              0.0 ns,
                              tperiod_WBLKB,
                              tpw_WBLKB_posedge,
                              tpw_WBLKB_negedge,
                              (TO_X01(WRB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9AST",
                              True,
                              True,
                              WARNING
                              );
 end if;

   ------------------------------------------------------------
   --               FIFO RESET                               --
   ------------------------------------------------------------

   if(RESET_ipd'event AND RESET_ipd = '0') then
       WADDR      := 0;
       RADDR      := 0;
       WADDR_wrap := 0;
       RADDR_wrap := 0;
       FULL_zd    := '0';
       EMPTY_tmp  := '1';
       EQTH_tmp   := '0';
       GEQTH_tmp  := '0';
       READ_AT_PREV_EDGE <='0';
       WPE_zd     := 'X';
       WB_initialized := False;
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
   end if;

   if ( RESET_ipd'event and RESET_ipd = '1' ) then
     if ( TO_X01 ( WBint ) = '0' ) then
       EMPTY_zd        := '0';
       EQTH_zd         := '1';
       GEQTH_zd        := '1';
       hold_empty_low  := 1;
       hold_eqth_high  := 1;
       hold_geqth_high := 1;
     end if;
   end if;

   if ( WBint'event ) then
     hold_empty_low  := 0;
     hold_eqth_high  := 0;
     hold_geqth_high := 0;
   end if;

   ------------------------------------------------------------
   --    wpe output                                           -
   ------------------------------------------------------------

   if ( PARODD_ipd'EVENT ) then
     WPE_zd   := not WPE_zd;
     RPE_zd   := not RPE_zd;
   end if;

   ------------------------------------------------------------
   --         WPE generating block                            -
   ------------------------------------------------------------

     tmp_par  := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;
     par_f  <= tmp_par ;
     tmp_par2 := (tmp_par xor DI8_ipd);
     par_f2  <=  tmp_par2;

     if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
         ( TO_X01 ( DI8_ipd )    = 'X' ) or
         ( TO_X01 ( DI7_ipd )    = 'X' ) or
         ( TO_X01 ( DI6_ipd )    = 'X' ) or
         ( TO_X01 ( DI5_ipd )    = 'X' ) or
         ( TO_X01 ( DI4_ipd )    = 'X' ) or
         ( TO_X01 ( DI3_ipd )    = 'X' ) or
         ( TO_X01 ( DI2_ipd )    = 'X' ) or
         ( TO_X01 ( DI1_ipd )    = 'X' ) or
         ( TO_X01 ( DI0_ipd )    = 'X' )
        ) then
       wpe_var  :=  'X';
     else
       if ( tmp_par2 /= PARODD_ipd ) then
         wpe_var  :=  '1';
       else
         wpe_var  :=  '0';
       end if;
     end if;
     RAM_di_int(8) := DI8_ipd;
     WPE_zd := wpe_var;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

   if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
   end if; 

   -----------------------------------------------------------
   --    calculate the depth and levels                     --
   -----------------------------------------------------------

    temp :=((INT(LGDEP2_delayed)*4) + (INT(LGDEP1_delayed)*2) + 
           (INT(LGDEP0_delayed)*1));

    case temp is 
         when 0 => depth := 2;
         when 1 => depth := 4;
         when 2 => depth := 8;
         when 3 => depth := 16;
         when 4 => depth := 32;
         when 5 => depth := 64;
         when 6 => depth := 128;
         when 7 => depth := 256;
         when others => depth := 0;
    end case;

    -- thresh value

    thresh := (INT(LEVEL7_delayed)*128) + (INT(LEVEL6_delayed)*64) + 
               (INT(LEVEL5_delayed)*32) + (INT(LEVEL4_delayed)*16) + 
               (INT(LEVEL3_delayed)*8) + (INT(LEVEL2_delayed)*4) + 
               (INT(LEVEL1_delayed)*2) + (INT(LEVEL0_delayed)*1); 

    if ( thresh = 0 or thresh = 255 ) then
      assert false
        report " Illegal level configuration, LEVEL cannot be 0 or 255 "
        severity failure;
    end if;

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

    if ( WBint'event AND WBint = '0') then
      if ( TO_X01 ( RESET_ipd ) = '1' ) then
        WB_initialized := True;
      end if;
    end if;

    if(WBint = '1') then
        null;
    elsif(WBint = '0') AND (TO_X01(RESET_ipd) = '1') then
        if(FULL_zd = '0') then 
        RAM_di_int(7 downto 0) := DI7_ipd & DI6_ipd & 
                                   DI5_ipd & DI4_ipd & 
                                   DI3_ipd & DI2_ipd & 
                                   DI1_ipd & DI0_ipd;
         memory_array(WADDR) := RAM_di_int;
       end if;
    else 
      null;
    end if;
    if (( WBint'event AND WBint = '1' ) AND 
        ( TO_X01 ( RESET_delayed ) = '1' ) AND
        ( WB_initialized )) then
      if(FULL_zd = '0') then 
       if(WADDR <depth-1  ) then
           WADDR := WADDR + 1;
       elsif( WADDR  = depth-1) then
         WADDR := 0;
         WADDR_wrap := 1 - WADDR_wrap;
       end if;
       if(WADDR   = RADDR ) then
         if(RADDR_wrap /= WADDR_wrap) then
            FULL_zd := '1';
            EMPTY_tmp :='0';
         end if;
       end if; 
         if(WADDR   /= RADDR ) then
          EMPTY_tmp := '0';
         end if;
          if(RADDR_wrap = WADDR_wrap) then
            if(WADDR - RADDR = thresh ) then
               EQTH_tmp := '1';
            else 
               EQTH_tmp := '0';
            end if;
            if(WADDR - RADDR >= thresh ) then
                GEQTH_tmp := '1';
            else 
                GEQTH_tmp := '0';
            end if;
          else 
           if((depth -RADDR + WADDR) = thresh ) then
               EQTH_tmp := '1';
           else 
               EQTH_tmp := '0';
           end if;
           if(depth - RADDR + WADDR >= thresh ) then
                GEQTH_tmp := '1';
           else 
                GEQTH_tmp := '0';
           end if;
         end if; 
        end if;
      end if;


  --------------------------------------------------------------------
  --          FIFO READ SECTION........                             --
  --------------------------------------------------------------------

  if (TO_X01(RCLKS_ipd)='X') then
    if(RESET_ipd /= '0') then
    if(TO_X01(RBint_delayed) /= '1') then
      if(TO_X01(RCLKS_previous) /= 'X') then
        assert false
        report ": RCLK unknown"
        severity Error;
        DO0_zd  := 'X';
        DO1_zd  := 'X';
        DO2_zd  := 'X';
        DO3_zd  := 'X';
        DO4_zd  := 'X';
        DO5_zd  := 'X';
        DO6_zd  := 'X';
        DO7_zd  := 'X';
        DO8_zd  := 'X';
      end if;
     end if;
    end if;
   elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='1') AND (TO_X01(RESET_delayed) = '1')) then
     READ_AT_PREV_EDGE <='0';
     case (TO_X01(RBint_delayed)) is
        when '1' =>
                null;
        when '0' =>
         if(TO_X01(EMPTY_zd) /= '1') then 
           DO0_zd  := memory_array(RADDR)(0);
           DO1_zd  := memory_array(RADDR)(1);
           DO2_zd  := memory_array(RADDR)(2);
           DO3_zd  := memory_array(RADDR)(3);
           DO4_zd  := memory_array(RADDR)(4);
           DO5_zd  := memory_array(RADDR)(5);
           DO6_zd  := memory_array(RADDR)(6);
           DO7_zd  := memory_array(RADDR)(7);
           DO8_zd  := memory_array(RADDR)(8);
           READ_AT_PREV_EDGE <='1';
           if(RADDR <depth-1  ) then
             RADDR := RADDR + 1;
           else
             RADDR :=(RADDR +1) mod  depth;
             RADDR_wrap :=1 - RADDR_wrap;
           end if;
            do_par  := DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR DO3_zd XOR
                       DO2_zd XOR DO1_zd XOR DO0_zd;
            par_f <= do_par;
            if (do_par = 'X') then
             RPE_zd := 'X';
            elsif (do_par /= PARODD_delayed) then
             RPE_zd  :=  '1';
            else
             RPE_zd  :=  '0';
            end if;
         end if;
     when others =>
       if (TO_X01(RBint_previous) /= 'X') then
        assert false
        report ": RDB or RBLKB unknown"
        severity Error;
        end if;
           DO0_zd  := 'X';
           DO1_zd  := 'X';
           DO2_zd  := 'X';
           DO3_zd  := 'X';
           DO4_zd  := 'X';
           DO5_zd  := 'X';
           DO6_zd  := 'X';
           DO7_zd  := 'X';
           DO8_zd  := 'X';
     end case;
  elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='0') AND (TO_X01(RESET_delayed) = '1') AND (TO_X01(READ_AT_PREV_EDGE) = '1')) then
   READ_AT_PREV_EDGE <='0';
   if(RADDR = WADDR ) then
    if(RADDR_wrap = WADDR_wrap) then
       EMPTY_tmp := '1';
       FULL_zd  := '0';
    end if;
   end if;
   if(RADDR /= WADDR ) then
    FULL_zd  := '0';
   end if;
    if(WADDR_wrap = RADDR_wrap ) then
     if((WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((WADDR - RADDR) >= thresh  ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    else 
     if((depth + WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((depth + WADDR - RADDR) >= thresh ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    end if;
 else 
    null;
 end if;

   -- Mimic odd silicon flag behavior coming out of RESET with WB low
   
   if ( hold_empty_low = 1 ) then
     EMPTY_zd := '0';
   else
     EMPTY_zd := EMPTY_tmp;
   end if;

   if ( hold_eqth_high = 1 ) then
     EQTH_zd := '1';
   else
     EQTH_zd := EQTH_tmp;
   end if;

   -- If LEVEL greater than DEPTH then GEQTH mimics FULL
   
   if ( hold_geqth_high = 1 ) then
     GEQTH_zd := '1';
   else
     if ( thresh > depth ) then
       GEQTH_zd := FULL_zd;
     else
       GEQTH_zd := GEQTH_tmp;
     end if;
   end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       RCLKS_previous   := RCLKS_ipd;
       RBint_previous   := RBint_delayed;
       RBint_delayed    := RBint;
       WBint_previous   := WBint;
       LGDEP0_previous  := LGDEP0_delayed;
       LGDEP0_delayed   := LGDEP0_ipd;
       LGDEP1_previous  := LGDEP1_delayed;
       LGDEP1_delayed   := LGDEP1_ipd;
       LGDEP2_previous  := LGDEP2_delayed;
       LGDEP2_delayed   := LGDEP2_ipd;
       LEVEL0_previous  := LEVEL0_delayed;
       LEVEL0_delayed   := LEVEL0_ipd;
       LEVEL1_previous  := LEVEL1_delayed;
       LEVEL1_delayed   := LEVEL1_ipd;
       LEVEL2_previous  := LEVEL2_delayed;
       LEVEL2_delayed   := LEVEL2_ipd;
       LEVEL3_previous  := LEVEL3_delayed;
       LEVEL3_delayed   := LEVEL3_ipd;
       LEVEL4_previous  := LEVEL4_delayed;
       LEVEL4_delayed   := LEVEL4_ipd;
       LEVEL5_previous  := LEVEL5_delayed;
       LEVEL5_delayed   := LEVEL5_ipd;
       LEVEL6_previous  := LEVEL6_delayed;
       LEVEL6_delayed   := LEVEL6_ipd;
       LEVEL7_previous  := LEVEL7_delayed;
       LEVEL7_delayed   := LEVEL7_ipd;
       PARODD_previous  := PARODD_delayed; 
       PARODD_delayed   := PARODD_ipd;
       RESET_previous   := RESET_delayed; 
       RESET_delayed    := RESET_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
             OutSignal     => DOS,
             GlitchData    => DOS_GlitchData,
             OutSignalName => "DOS",
             OutTemp       => DOS_zd,

             Paths =>   (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
           OutSignal     => WPE,
           GlitchData    => WPE_GlitchData,
           OutSignalName => "WPE",
           OutTemp       => WPE_zd,

           Paths =>   (0 => (DI0_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI0_WPE), true),
                       1 => (DI1_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI1_WPE), true),
                       2 => (DI2_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI2_WPE), true),
                       3 => (DI3_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI3_WPE), true),
                       4 => (DI4_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI4_WPE), true),
                       5 => (DI5_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI5_WPE), true),
                       6 => (DI6_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI6_WPE), true),
                       7 => (DI7_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI7_WPE), true),
                       8 => (DI8_ipd'last_event,
                                       VitalExtendToFillDelay(tpd_DI8_WPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO0), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO1), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO2), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO3), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO4), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO5), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO6), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO7), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO8), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => RPE,
           GlitchData    => RPE_GlitchData,
           OutSignalName => "RPE",
           OutTemp       => RPE_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_RPE), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_RPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => FULL,
           GlitchData    => FULL_GlitchData,
           OutSignalName => "FULL",
           OutTemp       => FULL_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_FULL), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_FULL), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_FULL), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_FULL), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EMPTY,
           GlitchData    => EMPTY_GlitchData,
           OutSignalName => "EMPTY",
           OutTemp       => EMPTY_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EMPTY), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_EMPTY), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_EMPTY), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EMPTY), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EQTH,
           GlitchData    => EQTH_GlitchData,
           OutSignalName => "EQTH",
           OutTemp       => EQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EQTH), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_EQTH), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_EQTH), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => GEQTH,
           GlitchData    => GEQTH_GlitchData,
           OutSignalName => "GEQTH",
           OutTemp       => GEQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_GEQTH), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_GEQTH), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_GEQTH), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_GEQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );


   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

LIBRARY a500k;
USE a500k.all;

entity FIFO256x9ASTP is 
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WRB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	thold_DI0_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI0_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI1_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI1_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI2_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI2_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI3_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI3_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI4_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI4_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI5_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI5_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI6_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI6_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI7_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI7_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI8_WRB_posedge_posedge                 : VitalDelayType := 0.000 ns;
	thold_DI8_WRB_negedge_posedge                 : VitalDelayType := 0.000 ns;
 	thold_DI0_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WBLKB_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WBLKB_negedge_posedge               : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI0_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI1_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI2_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI3_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI4_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI5_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI6_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI7_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WRB_posedge_posedge                : VitalDelayType := 0.000 ns;
	tsetup_DI8_WRB_negedge_posedge                : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WBLKB_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WBLKB_negedge_posedge              : VitalDelayType := 0.000 ns;

  	-- WB falling edge hold to RESETB   
 	thold_WRB_RESET_posedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_RESET_posedge_posedge             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_RESET_posedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_RESET_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_WRB_RESET_negedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WBLKB_RESET_negedge_posedge             : VitalDelayType := 0.000 ns;
	tsetup_WRB_RESET_negedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_RESET_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tpw_WRB_posedge                               : VitalDelayType := 0.000 ns;
 	tpw_WRB_negedge                               : VitalDelayType := 0.000 ns;
 	tperiod_WRB                                   : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WBLKB_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WBLKB                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');


ATTRIBUTE VITAL_LEVEL0 OF FIFO256x9ASTP : entity IS True ;
END FIFO256x9ASTP;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of FIFO256x9ASTP is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal LGDEP0_ipd : std_ulogic := 'X';
   signal LGDEP1_ipd : std_ulogic := 'X';
   signal LGDEP2_ipd : std_ulogic := 'X';
   signal LEVEL0_ipd : std_ulogic := 'X';
   signal LEVEL1_ipd : std_ulogic := 'X';
   signal LEVEL2_ipd : std_ulogic := 'X';
   signal LEVEL3_ipd : std_ulogic := 'X';
   signal LEVEL4_ipd : std_ulogic := 'X';
   signal LEVEL5_ipd : std_ulogic := 'X';
   signal LEVEL6_ipd : std_ulogic := 'X';
   signal LEVEL7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal RESET_ipd  : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

   -- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic := 'X';
   signal par_f2     : std_logic := 'X';

   signal WRITE_AT_PREV_EDGE : std_logic := '0';
   signal READ_AT_PREV_EDGE  : std_logic := '0';

   begin  --  VITAL_ACT

   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (LGDEP0_ipd, LGDEP0, VitalExtendToFillDelay(tipd_LGDEP0));
   VitalWireDelay (LGDEP1_ipd, LGDEP1, VitalExtendToFillDelay(tipd_LGDEP1));
   VitalWireDelay (LGDEP2_ipd, LGDEP2, VitalExtendToFillDelay(tipd_LGDEP2));
   VitalWireDelay (LEVEL0_ipd, LEVEL0, VitalExtendToFillDelay(tipd_LEVEL0));
   VitalWireDelay (LEVEL1_ipd, LEVEL1, VitalExtendToFillDelay(tipd_LEVEL1));
   VitalWireDelay (LEVEL2_ipd, LEVEL2, VitalExtendToFillDelay(tipd_LEVEL2));
   VitalWireDelay (LEVEL3_ipd, LEVEL3, VitalExtendToFillDelay(tipd_LEVEL3));
   VitalWireDelay (LEVEL4_ipd, LEVEL4, VitalExtendToFillDelay(tipd_LEVEL4));
   VitalWireDelay (LEVEL5_ipd, LEVEL5, VitalExtendToFillDelay(tipd_LEVEL5));
   VitalWireDelay (LEVEL6_ipd, LEVEL6, VitalExtendToFillDelay(tipd_LEVEL6));
   VitalWireDelay (LEVEL7_ipd, LEVEL7, VitalExtendToFillDelay(tipd_LEVEL7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RESET_ipd, RESET, VitalExtendToFillDelay(tipd_RESET));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

   ---------------------------------------------------------------
   --                  Behavior Section                         --
   ---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);

    VITALBehavior : process (
                          LEVEL0_ipd, LEVEL1_ipd, LEVEL2_ipd, LEVEL3_ipd, LEVEL4_ipd, LEVEL5_ipd, LEVEL6_ipd, LEVEL7_ipd, 
                          LGDEP0_ipd, LGDEP1_ipd, LGDEP2_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd, RESET_ipd
                          )

     -- some internal veriable declaration
     variable RAM_di_int   : std_logic_vector(8 downto 0);
     variable memory_array : MEM_TYPE  := (others =>(others => 'X'));
     variable do_par       : std_logic := 'X';
     variable tmp_par      : std_logic := 'X';
     variable tmp_par2     : std_logic := 'X';
     variable wpe_var      : std_logic := 'X';
     variable temp         : integer   := 0;
     variable thresh       : integer   := 0;
     variable depth        : integer   := 0;
     variable WADDR        : integer   := 0;
     variable WADDR_wrap   : integer   := 0;
     variable RADDR        : integer   := 0;
     variable RADDR_wrap   : integer   := 0;

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     --  Read Timing Check Results
     variable PeriodData_RESET           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET                : X01                 := '0';
     variable Tviol_PARODD_RCLKS_posedge : X01                 := '0';
     variable TmDt_PARODD_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_RCLKS_posedge  : X01                 := '0';
     variable Tmkr_RESET_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable PeriodData_WRB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WRB                  : X01                 := '0';
     variable PeriodData_WBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WBLKB                : X01                 := '0';
     variable Tviol_DI0_WRB_posedge      : X01                 := '0';
     variable TmDt_DI0_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI0_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI0_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WRB_posedge      : X01                 := '0';
     variable TmDt_DI1_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI1_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WRB_posedge      : X01                 := '0';
     variable TmDt_DI2_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI2_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WRB_posedge      : X01                 := '0';
     variable TmDt_DI3_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI3_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WRB_posedge      : X01                 := '0';
     variable TmDt_DI4_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI4_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WRB_posedge      : X01                 := '0';
     variable TmDt_DI5_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI5_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WRB_posedge      : X01                 := '0';
     variable TmDt_DI6_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI6_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WRB_posedge      : X01                 := '0';
     variable TmDt_DI7_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI7_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WRB_posedge      : X01                 := '0';
     variable TmDt_DI8_WRB_posedge       : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WBLKB_posedge    : X01                 := '0';
     variable TmDt_DI8_WBLKB_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_RESET_posedge    : X01                 := '0';
     variable TmDt_WRB_RESET_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_RESET_posedge  : X01                 := '0';
     variable TmDt_WBLKB_RESET_posedge   : VitalTimingDataType := VitalTimingDataInit;

     -- functional Results


     variable DO0_zd   : std_ulogic;
     variable DO1_zd   : std_ulogic;
     variable DO2_zd   : std_ulogic;
     variable DO3_zd   : std_ulogic;
     variable DO4_zd   : std_ulogic;
     variable DO5_zd   : std_ulogic;
     variable DO6_zd   : std_ulogic;
     variable DO7_zd   : std_ulogic;
     variable DO8_zd   : std_ulogic;
     variable RPE_zd   : std_ulogic;
     variable WPE_zd   : std_ulogic;
     variable DOS_zd   : std_ulogic;
     variable FULL_zd  : std_ulogic;
     variable EMPTY_zd : std_ulogic;
     variable EQTH_zd  : std_ulogic;
     variable GEQTH_zd : std_ulogic;
     variable EMPTY_tmp : std_ulogic;
     variable EQTH_tmp  : std_ulogic;
     variable GEQTH_tmp : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData   : VitalGlitchDataType;
     variable DO1_GlitchData   : VitalGlitchDataType;
     variable DO2_GlitchData   : VitalGlitchDataType;
     variable DO3_GlitchData   : VitalGlitchDataType;
     variable DO4_GlitchData   : VitalGlitchDataType;
     variable DO5_GlitchData   : VitalGlitchDataType;
     variable DO6_GlitchData   : VitalGlitchDataType;
     variable DO7_GlitchData   : VitalGlitchDataType;
     variable DO8_GlitchData   : VitalGlitchDataType;
     variable DOS_GlitchData   : VitalGlitchDataType;
     variable FULL_GlitchData  : VitalGlitchDataType;
     variable EMPTY_GlitchData : VitalGlitchDataType;
     variable EQTH_GlitchData  : VitalGlitchDataType;
     variable GEQTH_GlitchData : VitalGlitchDataType;

     -- last value variables
     variable RCLKS_previous   : std_ulogic := 'X';
     variable RBint_delayed    : std_ulogic := 'X';
     variable RBint_previous   : std_ulogic := 'X';
     variable WBint_previous   : std_ulogic := 'X';
     variable DIS_previous     : std_ulogic := 'X';
     variable RESET_previous   : std_ulogic := 'X';
     variable RESET_delayed    : std_ulogic := 'X';
     variable PARODD_previous  : std_ulogic := 'X';
     variable PARODD_delayed   : std_ulogic := 'X';
     variable DI0_delayed      : std_ulogic := 'X';
     variable DI1_delayed      : std_ulogic := 'X';
     variable DI2_delayed      : std_ulogic := 'X';
     variable DI3_delayed      : std_ulogic := 'X';
     variable DI4_delayed      : std_ulogic := 'X';
     variable DI5_delayed      : std_ulogic := 'X';
     variable DI6_delayed      : std_ulogic := 'X';
     variable DI7_delayed      : std_ulogic := 'X';
     variable DI8_delayed      : std_ulogic := 'X';
     variable DI0_previous     : std_ulogic := 'X';
     variable DI1_previous     : std_ulogic := 'X';
     variable DI2_previous     : std_ulogic := 'X';
     variable DI3_previous     : std_ulogic := 'X';
     variable DI4_previous     : std_ulogic := 'X';
     variable DI5_previous     : std_ulogic := 'X';
     variable DI6_previous     : std_ulogic := 'X';
     variable DI7_previous     : std_ulogic := 'X';
     variable DI8_previous     : std_ulogic := 'X';
     variable LGDEP0_delayed   : std_ulogic := 'X';
     variable LGDEP1_delayed   : std_ulogic := 'X';
     variable LGDEP2_delayed   : std_ulogic := 'X';
     variable LGDEP0_previous  : std_ulogic := 'X';
     variable LGDEP1_previous  : std_ulogic := 'X';
     variable LGDEP2_previous  : std_ulogic := 'X';
     variable LEVEL0_delayed   : std_ulogic := 'X';
     variable LEVEL1_delayed   : std_ulogic := 'X';
     variable LEVEL2_delayed   : std_ulogic := 'X';
     variable LEVEL3_delayed   : std_ulogic := 'X';
     variable LEVEL4_delayed   : std_ulogic := 'X';
     variable LEVEL5_delayed   : std_ulogic := 'X';
     variable LEVEL6_delayed   : std_ulogic := 'X';
     variable LEVEL7_delayed   : std_ulogic := 'X';
     variable LEVEL0_previous  : std_ulogic := 'X';
     variable LEVEL1_previous  : std_ulogic := 'X';
     variable LEVEL2_previous  : std_ulogic := 'X';
     variable LEVEL3_previous  : std_ulogic := 'X';
     variable LEVEL4_previous  : std_ulogic := 'X';
     variable LEVEL5_previous  : std_ulogic := 'X';
     variable LEVEL6_previous  : std_ulogic := 'X';
     variable LEVEL7_previous  : std_ulogic := 'X';

     variable WB_initialized   : Boolean := False; 
     -- True = WB_int falling edge occured.  
     -- Must occur before first write after RESET.

     -- Special variables to control flags
     variable hold_empty_low   : integer := 0;
     variable hold_eqth_high   : integer := 0;
     variable hold_geqth_high  : integer := 0;

 begin -- process VITALBehavior

 if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

   -- recovery / removal check for RCLKS to RESET signal ;
       VitalRecoveryRemovalCheck ( Tviol_RESET_RCLKS_posedge,
                             Tmkr_RESET_RCLKS_posedge,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             trecovery_RESET_RCLKS_posedge_negedge,
                             thold_RESET_RCLKS_posedge_posedge,
                             TRUE,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'), 
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             TRUE,
                             TRUE,
                             WARNING
                             );

   -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             ((TO_X01(RBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             ((TO_X01(RDB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_PARODD_RCLKS_posedge,
                             TmDt_PARODD_RCLKS_posedge,
                             PARODD_ipd, "PARODD",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_PARODD_RCLKS_posedge_posedge,
                             tsetup_PARODD_RCLKS_negedge_posedge,
                             thold_PARODD_RCLKS_posedge_posedge,
                             thold_PARODD_RCLKS_negedge_posedge,
                             (TO_X01(RESET_ipd) = '1'),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (TO_X01(RDB) = '0') AND (TO_X01(RBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9ASTP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RESET,
                              PeriodData_RESET,
                              RESET_ipd, "RESET",
                              0.0 ns,
                              tpw_RESET_negedge,
                              0.0 ns,
                              tpw_RESET_negedge,
                              True,
                              InstancePath & "/FIFO256x9ASTP",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

   -- setup /hold check for WRB/WBLKB to RESET signal ;
       VitalSetupHoldCheck ( Tviol_WRB_RESET_posedge,
                             TmDt_WRB_RESET_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             tsetup_WRB_RESET_posedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             thold_WRB_RESET_negedge_posedge,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_RESET_posedge,
                             TmDt_WBLKB_RESET_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             tsetup_WBLKB_RESET_posedge_posedge,
                             0.0 ns,
                             0.0 ns,
                             thold_WBLKB_RESET_negedge_posedge,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WRB_posedge,
                             TmDt_DI0_WRB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI0_WRB_posedge_posedge,
                             tsetup_DI0_WRB_negedge_posedge,
                             thold_DI0_WRB_posedge_posedge,
                             thold_DI0_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WRB_posedge,
                             TmDt_DI1_WRB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI1_WRB_posedge_posedge,
                             tsetup_DI1_WRB_negedge_posedge,
                             thold_DI1_WRB_posedge_posedge,
                             thold_DI1_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WRB_posedge,
                             TmDt_DI2_WRB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI2_WRB_posedge_posedge,
                             tsetup_DI2_WRB_negedge_posedge,
                             thold_DI2_WRB_posedge_posedge,
                             thold_DI2_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WRB_posedge,
                             TmDt_DI3_WRB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI3_WRB_posedge_posedge,
                             tsetup_DI3_WRB_negedge_posedge,
                             thold_DI3_WRB_posedge_posedge,
                             thold_DI3_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WRB_posedge,
                             TmDt_DI4_WRB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI4_WRB_posedge_posedge,
                             tsetup_DI4_WRB_negedge_posedge,
                             thold_DI4_WRB_posedge_posedge,
                             thold_DI4_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WRB_posedge,
                             TmDt_DI5_WRB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI5_WRB_posedge_posedge,
                             tsetup_DI5_WRB_negedge_posedge,
                             thold_DI5_WRB_posedge_posedge,
                             thold_DI5_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WRB_posedge,
                             TmDt_DI6_WRB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI6_WRB_posedge_posedge,
                             tsetup_DI6_WRB_negedge_posedge,
                             thold_DI6_WRB_posedge_posedge,
                             thold_DI6_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WRB_posedge,
                             TmDt_DI7_WRB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI7_WRB_posedge_posedge,
                             tsetup_DI7_WRB_negedge_posedge,
                             thold_DI7_WRB_posedge_posedge,
                             thold_DI7_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WRB_posedge,
                             TmDt_DI8_WRB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WRB_ipd, "WRB",
                             0.0 ns, 
                             tsetup_DI8_WRB_posedge_posedge,
                             tsetup_DI8_WRB_negedge_posedge,
                             thold_DI8_WRB_posedge_posedge,
                             thold_DI8_WRB_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WBLKB_posedge,
                             TmDt_DI0_WBLKB_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI0_WBLKB_posedge_posedge,
                             tsetup_DI0_WBLKB_negedge_posedge,
                             thold_DI0_WBLKB_posedge_posedge,
                             thold_DI0_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI1_WBLKB_posedge,
                             TmDt_DI1_WBLKB_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI1_WBLKB_posedge_posedge,
                             tsetup_DI1_WBLKB_negedge_posedge,
                             thold_DI1_WBLKB_posedge_posedge,
                             thold_DI1_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI2_WBLKB_posedge,
                             TmDt_DI2_WBLKB_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI2_WBLKB_posedge_posedge,
                             tsetup_DI2_WBLKB_negedge_posedge,
                             thold_DI2_WBLKB_posedge_posedge,
                             thold_DI2_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI3_WBLKB_posedge,
                             TmDt_DI3_WBLKB_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI3_WBLKB_posedge_posedge,
                             tsetup_DI3_WBLKB_negedge_posedge,
                             thold_DI3_WBLKB_posedge_posedge,
                             thold_DI3_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI4_WBLKB_posedge,
                             TmDt_DI4_WBLKB_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI4_WBLKB_posedge_posedge,
                             tsetup_DI4_WBLKB_negedge_posedge,
                             thold_DI4_WBLKB_posedge_posedge,
                             thold_DI4_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI5_WBLKB_posedge,
                             TmDt_DI5_WBLKB_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI5_WBLKB_posedge_posedge,
                             tsetup_DI5_WBLKB_negedge_posedge,
                             thold_DI5_WBLKB_posedge_posedge,
                             thold_DI5_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI6_WBLKB_posedge,
                             TmDt_DI6_WBLKB_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI6_WBLKB_posedge_posedge,
                             tsetup_DI6_WBLKB_negedge_posedge,
                             thold_DI6_WBLKB_posedge_posedge,
                             thold_DI6_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI7_WBLKB_posedge,
                             TmDt_DI7_WBLKB_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI7_WBLKB_posedge_posedge,
                             tsetup_DI7_WBLKB_negedge_posedge,
                             thold_DI7_WBLKB_posedge_posedge,
                             thold_DI7_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
       VitalSetupHoldCheck ( Tviol_DI8_WBLKB_posedge,
                             TmDt_DI8_WBLKB_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns, 
                             tsetup_DI8_WBLKB_posedge_posedge,
                             tsetup_DI8_WBLKB_negedge_posedge,
                             thold_DI8_WBLKB_posedge_posedge,
                             thold_DI8_WBLKB_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9ASTP",
                             True,
                             True,
                             WARNING
                             );
      VitalPeriodPulseCheck ( Pviol_WRB,
                              PeriodData_WRB,
                              WRB_ipd, "WRB",
                              0.0 ns,
                              tperiod_WRB,
                              tpw_WRB_posedge,
                              tpw_WRB_negedge,
                              (TO_X01(WBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9ASTP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_WBLKB,
                              PeriodData_WBLKB,
                              WBLKB_ipd, "WBLKB",
                              0.0 ns,
                              tperiod_WBLKB,
                              tpw_WBLKB_posedge,
                              tpw_WBLKB_negedge,
                              (TO_X01(WRB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9ASTP",
                              True,
                              True,
                              WARNING
                              );
 end if;

   ------------------------------------------------------------
   --               FIFO RESET                               --
   ------------------------------------------------------------

   if(RESET_ipd'event AND RESET_ipd = '0') then
       WADDR      := 0;
       RADDR      := 0;
       WADDR_wrap := 0;
       RADDR_wrap := 0;
       FULL_zd    := '0';
       EMPTY_tmp  := '1';
       EQTH_tmp   := '0';
       GEQTH_tmp  := '0';
       READ_AT_PREV_EDGE <='0';
       WB_initialized := False;
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
   end if;

   if ( RESET_ipd'event and RESET_ipd = '1' ) then
     if ( TO_X01 ( WBint ) = '0' ) then
       EMPTY_zd        := '0';
       EQTH_zd         := '1';
       GEQTH_zd        := '1';
       hold_empty_low  := 1;
       hold_eqth_high  := 1;
       hold_geqth_high := 1;
     end if;
   end if;

   if ( WBint'event ) then
     hold_empty_low  := 0;
     hold_eqth_high  := 0;
     hold_geqth_high := 0;
   end if;

   ------------------------------------------------------------
   --         WPE generating block                            -
   ------------------------------------------------------------

     tmp_par  := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;
     par_f  <= tmp_par ;
     if (tmp_par /= PARODD_ipd) then
        wpe_var  :=  '1';
     else
        wpe_var  :=  '0';
     end if;
     RAM_di_int(8) := wpe_var;
     WPE_zd := wpe_var;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

   if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
   end if; 

   -----------------------------------------------------------
   --    calculate the depth and levels                     --
   -----------------------------------------------------------

    temp :=((INT(LGDEP2_delayed)*4) + (INT(LGDEP1_delayed)*2) + 
           (INT(LGDEP0_delayed)*1));

    case temp is 
         when 0 => depth := 2;
         when 1 => depth := 4;
         when 2 => depth := 8;
         when 3 => depth := 16;
         when 4 => depth := 32;
         when 5 => depth := 64;
         when 6 => depth := 128;
         when 7 => depth := 256;
         when others => depth := 0;
    end case;

    -- thresh value

    thresh := (INT(LEVEL7_delayed)*128) + (INT(LEVEL6_delayed)*64) + 
               (INT(LEVEL5_delayed)*32) + (INT(LEVEL4_delayed)*16) + 
               (INT(LEVEL3_delayed)*8) + (INT(LEVEL2_delayed)*4) + 
               (INT(LEVEL1_delayed)*2) + (INT(LEVEL0_delayed)*1); 

    if ( thresh = 0 or thresh = 255 ) then
      assert false
        report " Illegal level configuration, LEVEL cannot be 0 or 255 "
        severity failure;
    end if;

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

    if ( WBint'event AND WBint = '0') then
      if ( TO_X01 ( RESET_ipd ) = '1' ) then
        WB_initialized := True;
      end if;
    end if;

    if(WBint = '1') then
        null;
    elsif(WBint = '0') AND (TO_X01(RESET_ipd) = '1') then
        if(FULL_zd = '0') then 
        RAM_di_int(7 downto 0) := DI7_ipd & DI6_ipd & 
                                   DI5_ipd & DI4_ipd & 
                                   DI3_ipd & DI2_ipd & 
                                   DI1_ipd & DI0_ipd;
         memory_array(WADDR) := RAM_di_int;
       end if;
    else 
      null;
    end if;
    if (( WBint'event AND WBint = '1' ) AND 
        ( TO_X01 ( RESET_delayed ) = '1' ) AND
        ( WB_initialized )) then
      if(FULL_zd = '0') then 
       if(WADDR <depth-1  ) then
           WADDR := WADDR + 1;
       elsif( WADDR  = depth-1) then
         WADDR := 0;
         WADDR_wrap := 1 - WADDR_wrap;
       end if;
       if(WADDR   = RADDR ) then
         if(RADDR_wrap /= WADDR_wrap) then
            FULL_zd := '1';
            EMPTY_tmp :='0';
         end if;
       end if; 
         if(WADDR   /= RADDR ) then
          EMPTY_tmp := '0';
         end if;
          if(RADDR_wrap = WADDR_wrap) then
            if(WADDR - RADDR = thresh ) then
               EQTH_tmp := '1';
            else 
               EQTH_tmp := '0';
            end if;
            if(WADDR - RADDR >= thresh ) then
                GEQTH_tmp := '1';
            else 
                GEQTH_tmp := '0';
            end if;
          else 
           if((depth -RADDR + WADDR) = thresh ) then
               EQTH_tmp := '1';
           else 
               EQTH_tmp := '0';
           end if;
           if(depth - RADDR + WADDR >= thresh ) then
                GEQTH_tmp := '1';
           else 
                GEQTH_tmp := '0';
           end if;
         end if; 
        end if;
      end if;


  --------------------------------------------------------------------
  --          FIFO READ SECTION........                             --
  --------------------------------------------------------------------

  if (TO_X01(RCLKS_ipd)='X') then
    if(RESET_ipd /= '0') then
    if(TO_X01(RBint_delayed) /= '1') then
      if(TO_X01(RCLKS_previous) /= 'X') then
        assert false
        report ": RCLK unknown"
        severity Error;
        DO0_zd  := 'X';
        DO1_zd  := 'X';
        DO2_zd  := 'X';
        DO3_zd  := 'X';
        DO4_zd  := 'X';
        DO5_zd  := 'X';
        DO6_zd  := 'X';
        DO7_zd  := 'X';
        DO8_zd  := 'X';
      end if;
     end if;
    end if;
   elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='1') AND (TO_X01(RESET_delayed) = '1')) then
     READ_AT_PREV_EDGE <='0';
     case (TO_X01(RBint_delayed)) is
        when '1' =>
                null;
        when '0' =>
         if(TO_X01(EMPTY_zd) /= '1') then 
           DO0_zd  := memory_array(RADDR)(0);
           DO1_zd  := memory_array(RADDR)(1);
           DO2_zd  := memory_array(RADDR)(2);
           DO3_zd  := memory_array(RADDR)(3);
           DO4_zd  := memory_array(RADDR)(4);
           DO5_zd  := memory_array(RADDR)(5);
           DO6_zd  := memory_array(RADDR)(6);
           DO7_zd  := memory_array(RADDR)(7);
           DO8_zd  := memory_array(RADDR)(8);
           READ_AT_PREV_EDGE <='1';
           if(RADDR <depth-1  ) then
             RADDR := RADDR + 1;
           else
             RADDR :=(RADDR +1) mod  depth;
             RADDR_wrap :=1 - RADDR_wrap;
           end if;
            do_par  := DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR DO3_zd XOR
                       DO2_zd XOR DO1_zd XOR DO0_zd;
            par_f <= do_par;
            if (do_par = 'X') then
             RPE_zd := 'X';
            elsif (do_par /= PARODD_delayed) then
             RPE_zd  :=  '1';
            else
             RPE_zd  :=  '0';
            end if;
         end if;
     when others =>
       if (TO_X01(RBint_previous) /= 'X') then
        assert false
        report ": RDB or RBLKB unknown"
        severity Error;
        end if;
           DO0_zd  := 'X';
           DO1_zd  := 'X';
           DO2_zd  := 'X';
           DO3_zd  := 'X';
           DO4_zd  := 'X';
           DO5_zd  := 'X';
           DO6_zd  := 'X';
           DO7_zd  := 'X';
           DO8_zd  := 'X';
     end case;
  elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='0') AND (TO_X01(RESET_delayed) = '1') AND (TO_X01(READ_AT_PREV_EDGE) = '1')) then
   READ_AT_PREV_EDGE <='0';
   if(RADDR = WADDR ) then
    if(RADDR_wrap = WADDR_wrap) then
       EMPTY_tmp := '1';
       FULL_zd  := '0';
    end if;
   end if;
   if(RADDR /= WADDR ) then
    FULL_zd  := '0';
   end if;
    if(WADDR_wrap = RADDR_wrap ) then
     if((WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((WADDR - RADDR) >= thresh  ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    else 
     if((depth + WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((depth + WADDR - RADDR) >= thresh ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    end if;
 else 
    null;
 end if;


   -- Mimic odd silicon flag behavior coming out of RESET with WB low
   
   if ( hold_empty_low = 1 ) then
     EMPTY_zd := '0';
   else
     EMPTY_zd := EMPTY_tmp;
   end if;

   if ( hold_eqth_high = 1 ) then
     EQTH_zd := '1';
   else
     EQTH_zd := EQTH_tmp;
   end if;

   -- If LEVEL greater than DEPTH then GEQTH mimics FULL
   
   if ( hold_geqth_high = 1 ) then
     GEQTH_zd := '1';
   else
     if ( thresh > depth ) then
       GEQTH_zd := FULL_zd;
     else
       GEQTH_zd := GEQTH_tmp;
     end if;
   end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       RCLKS_previous   := RCLKS_ipd;
       RBint_previous   := RBint_delayed;
       RBint_delayed    := RBint;
       WBint_previous   := WBint;
       LGDEP0_previous  := LGDEP0_delayed;
       LGDEP0_delayed   := LGDEP0_ipd;
       LGDEP1_previous  := LGDEP1_delayed;
       LGDEP1_delayed   := LGDEP1_ipd;
       LGDEP2_previous  := LGDEP2_delayed;
       LGDEP2_delayed   := LGDEP2_ipd;
       LEVEL0_previous  := LEVEL0_delayed;
       LEVEL0_delayed   := LEVEL0_ipd;
       LEVEL1_previous  := LEVEL1_delayed;
       LEVEL1_delayed   := LEVEL1_ipd;
       LEVEL2_previous  := LEVEL2_delayed;
       LEVEL2_delayed   := LEVEL2_ipd;
       LEVEL3_previous  := LEVEL3_delayed;
       LEVEL3_delayed   := LEVEL3_ipd;
       LEVEL4_previous  := LEVEL4_delayed;
       LEVEL4_delayed   := LEVEL4_ipd;
       LEVEL5_previous  := LEVEL5_delayed;
       LEVEL5_delayed   := LEVEL5_ipd;
       LEVEL6_previous  := LEVEL6_delayed;
       LEVEL6_delayed   := LEVEL6_ipd;
       LEVEL7_previous  := LEVEL7_delayed;
       LEVEL7_delayed   := LEVEL7_ipd;
       PARODD_previous  := PARODD_delayed; 
       PARODD_delayed   := PARODD_ipd;
       RESET_previous   := RESET_delayed; 
       RESET_delayed    := RESET_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
             OutSignal     => DOS,
             GlitchData    => DOS_GlitchData,
             OutSignalName => "DOS",
             OutTemp       => DOS_zd,

             Paths =>   (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO0), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO1), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO2), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO3), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO4), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO5), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO6), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO7), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO8), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => FULL,
           GlitchData    => FULL_GlitchData,
           OutSignalName => "FULL",
           OutTemp       => FULL_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_FULL), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_FULL), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_FULL), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_FULL), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EMPTY,
           GlitchData    => EMPTY_GlitchData,
           OutSignalName => "EMPTY",
           OutTemp       => EMPTY_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EMPTY), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_EMPTY), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_EMPTY), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EMPTY), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EQTH,
           GlitchData    => EQTH_GlitchData,
           OutSignalName => "EQTH",
           OutTemp       => EQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EQTH), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_EQTH), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_EQTH), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => GEQTH,
           GlitchData    => GEQTH_GlitchData,
           OutSignalName => "GEQTH",
           OutTemp       => GEQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_GEQTH), true),
                       1 => (WRB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WRB_GEQTH), true),
                       2 => (WBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WBLKB_GEQTH), true),
                       3 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_GEQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );


   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

LIBRARY a500k;
USE a500k.all;

entity FIFO256x9SA is 
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_PARODD_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tpw_RDB_posedge         : VitalDelayType        := 0.000 ns;
 	tpw_RDB_negedge         : VitalDelayType        := 0.000 ns;
 	tperiod_RDB             : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_posedge       : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_negedge       : VitalDelayType        := 0.000 ns;
 	tperiod_RBLKB           : VitalDelayType        := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_WCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_WCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;

        -- WCLK falling edge setup to RESET rising edge 
 	trecovery_RESET_WCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_WCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- WCLK rising  edge hold to RESET rising edge 
	thold_RESET_WCLKS_posedge_posedge             : VitalDelayType := 0.00 ns;
	thold_RESET_WCLKS_posedge_negedge             : VitalDelayType := 0.00 ns;
	tpw_WCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        WPE    :  OUT STD_LOGIC := 'X';
        RPE    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        WCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');


ATTRIBUTE VITAL_LEVEL0 OF FIFO256x9SA : entity IS True ;
END FIFO256x9SA;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of FIFO256x9SA is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal LGDEP0_ipd : std_ulogic := 'X';
   signal LGDEP1_ipd : std_ulogic := 'X';
   signal LGDEP2_ipd : std_ulogic := 'X';
   signal LEVEL0_ipd : std_ulogic := 'X';
   signal LEVEL1_ipd : std_ulogic := 'X';
   signal LEVEL2_ipd : std_ulogic := 'X';
   signal LEVEL3_ipd : std_ulogic := 'X';
   signal LEVEL4_ipd : std_ulogic := 'X';
   signal LEVEL5_ipd : std_ulogic := 'X';
   signal LEVEL6_ipd : std_ulogic := 'X';
   signal LEVEL7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal RESET_ipd  : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal WCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

   -- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic := 'X';
   signal par_f2     : std_logic := 'X';

   signal WRITE_AT_PREV_EDGE : std_logic := '0';
   signal READ_AT_PREV_EDGE  : std_logic := '0';

   begin  --  VITAL_ACT

   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (LGDEP0_ipd, LGDEP0, VitalExtendToFillDelay(tipd_LGDEP0));
   VitalWireDelay (LGDEP1_ipd, LGDEP1, VitalExtendToFillDelay(tipd_LGDEP1));
   VitalWireDelay (LGDEP2_ipd, LGDEP2, VitalExtendToFillDelay(tipd_LGDEP2));
   VitalWireDelay (LEVEL0_ipd, LEVEL0, VitalExtendToFillDelay(tipd_LEVEL0));
   VitalWireDelay (LEVEL1_ipd, LEVEL1, VitalExtendToFillDelay(tipd_LEVEL1));
   VitalWireDelay (LEVEL2_ipd, LEVEL2, VitalExtendToFillDelay(tipd_LEVEL2));
   VitalWireDelay (LEVEL3_ipd, LEVEL3, VitalExtendToFillDelay(tipd_LEVEL3));
   VitalWireDelay (LEVEL4_ipd, LEVEL4, VitalExtendToFillDelay(tipd_LEVEL4));
   VitalWireDelay (LEVEL5_ipd, LEVEL5, VitalExtendToFillDelay(tipd_LEVEL5));
   VitalWireDelay (LEVEL6_ipd, LEVEL6, VitalExtendToFillDelay(tipd_LEVEL6));
   VitalWireDelay (LEVEL7_ipd, LEVEL7, VitalExtendToFillDelay(tipd_LEVEL7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RESET_ipd, RESET, VitalExtendToFillDelay(tipd_RESET));
   VitalWireDelay (WCLKS_ipd, WCLKS, VitalExtendToFillDelay(tipd_WCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

   ---------------------------------------------------------------
   --                  Behavior Section                         --
   ---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);

    VITALBehavior : process (
                          LEVEL0_ipd, LEVEL1_ipd, LEVEL2_ipd, LEVEL3_ipd, LEVEL4_ipd, LEVEL5_ipd, LEVEL6_ipd, LEVEL7_ipd, 
                          LGDEP0_ipd, LGDEP1_ipd, LGDEP2_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          WCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd, RESET_ipd
                          )

     -- some internal veriable declaration
     variable RAM_di_int   : std_logic_vector(8 downto 0);
     variable memory_array : MEM_TYPE  := (others =>(others => 'X'));
     variable do_par       : std_logic := 'X';
     variable tmp_par      : std_logic := 'X';
     variable tmp_par2     : std_logic := 'X';
     variable wpe_var      : std_logic := 'X';
     variable temp         : integer   := 0;
     variable thresh       : integer   := 0;
     variable depth        : integer   := 0;
     variable WADDR        : integer   := 0;
     variable WADDR_wrap   : integer   := 0;
     variable RADDR        : integer   := 0;
     variable RADDR_wrap   : integer   := 0;

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     --  Read Timing Check Results
     variable PeriodData_RESET           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET                : X01                 := '0';
     variable PeriodData_RDB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RDB                  : X01                 := '0';
     variable PeriodData_RBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RBLKB                : X01                 := '0';
     variable Tviol_DI0_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI0_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI1_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI2_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI3_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI4_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI5_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI6_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI7_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI8_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_PARODD_WCLKS_posedge : X01                 := '0';
     variable TmDt_PARODD_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_WCLKS_posedge    : X01                 := '0';
     variable TmDt_WRB_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_WCLKS_posedge  : X01                 := '0';
     variable TmDt_WBLKB_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_WCLKS_posedge  : X01                 := '0';
     variable Tmkr_RESET_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WCLKS                : X01                 := '0';

     -- functional Results


     variable DO0_zd   : std_ulogic;
     variable DO1_zd   : std_ulogic;
     variable DO2_zd   : std_ulogic;
     variable DO3_zd   : std_ulogic;
     variable DO4_zd   : std_ulogic;
     variable DO5_zd   : std_ulogic;
     variable DO6_zd   : std_ulogic;
     variable DO7_zd   : std_ulogic;
     variable DO8_zd   : std_ulogic;
     variable RPE_zd   : std_ulogic;
     variable WPE_zd   : std_ulogic;
     variable DOS_zd   : std_ulogic;
     variable FULL_zd  : std_ulogic;
     variable EMPTY_zd : std_ulogic;
     variable EQTH_zd  : std_ulogic;
     variable GEQTH_zd : std_ulogic;
     variable FULL_tmp  : std_ulogic;
     variable EMPTY_tmp : std_ulogic;
     variable EQTH_tmp  : std_ulogic;
     variable GEQTH_tmp : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData   : VitalGlitchDataType;
     variable DO1_GlitchData   : VitalGlitchDataType;
     variable DO2_GlitchData   : VitalGlitchDataType;
     variable DO3_GlitchData   : VitalGlitchDataType;
     variable DO4_GlitchData   : VitalGlitchDataType;
     variable DO5_GlitchData   : VitalGlitchDataType;
     variable DO6_GlitchData   : VitalGlitchDataType;
     variable DO7_GlitchData   : VitalGlitchDataType;
     variable DO8_GlitchData   : VitalGlitchDataType;
     variable RPE_GlitchData   : VitalGlitchDataType;
     variable WPE_GlitchData   : VitalGlitchDataType;
     variable DOS_GlitchData   : VitalGlitchDataType;
     variable FULL_GlitchData  : VitalGlitchDataType;
     variable EMPTY_GlitchData : VitalGlitchDataType;
     variable EQTH_GlitchData  : VitalGlitchDataType;
     variable GEQTH_GlitchData : VitalGlitchDataType;

     -- last value variables
     variable WCLKS_previous   : std_ulogic := 'X';
     variable RBint_previous   : std_ulogic := 'X';
     variable WBint_delayed    : std_ulogic := 'X';
     variable WBint_previous   : std_ulogic := 'X';
     variable DIS_previous     : std_ulogic := 'X';
     variable RESET_previous   : std_ulogic := 'X';
     variable RESET_delayed    : std_ulogic := 'X';
     variable PARODD_previous  : std_ulogic := 'X';
     variable PARODD_delayed   : std_ulogic := 'X';
     variable DI0_delayed      : std_ulogic := 'X';
     variable DI1_delayed      : std_ulogic := 'X';
     variable DI2_delayed      : std_ulogic := 'X';
     variable DI3_delayed      : std_ulogic := 'X';
     variable DI4_delayed      : std_ulogic := 'X';
     variable DI5_delayed      : std_ulogic := 'X';
     variable DI6_delayed      : std_ulogic := 'X';
     variable DI7_delayed      : std_ulogic := 'X';
     variable DI8_delayed      : std_ulogic := 'X';
     variable DI0_previous     : std_ulogic := 'X';
     variable DI1_previous     : std_ulogic := 'X';
     variable DI2_previous     : std_ulogic := 'X';
     variable DI3_previous     : std_ulogic := 'X';
     variable DI4_previous     : std_ulogic := 'X';
     variable DI5_previous     : std_ulogic := 'X';
     variable DI6_previous     : std_ulogic := 'X';
     variable DI7_previous     : std_ulogic := 'X';
     variable DI8_previous     : std_ulogic := 'X';
     variable LGDEP0_delayed   : std_ulogic := 'X';
     variable LGDEP1_delayed   : std_ulogic := 'X';
     variable LGDEP2_delayed   : std_ulogic := 'X';
     variable LGDEP0_previous  : std_ulogic := 'X';
     variable LGDEP1_previous  : std_ulogic := 'X';
     variable LGDEP2_previous  : std_ulogic := 'X';
     variable LEVEL0_delayed   : std_ulogic := 'X';
     variable LEVEL1_delayed   : std_ulogic := 'X';
     variable LEVEL2_delayed   : std_ulogic := 'X';
     variable LEVEL3_delayed   : std_ulogic := 'X';
     variable LEVEL4_delayed   : std_ulogic := 'X';
     variable LEVEL5_delayed   : std_ulogic := 'X';
     variable LEVEL6_delayed   : std_ulogic := 'X';
     variable LEVEL7_delayed   : std_ulogic := 'X';
     variable LEVEL0_previous  : std_ulogic := 'X';
     variable LEVEL1_previous  : std_ulogic := 'X';
     variable LEVEL2_previous  : std_ulogic := 'X';
     variable LEVEL3_previous  : std_ulogic := 'X';
     variable LEVEL4_previous  : std_ulogic := 'X';
     variable LEVEL5_previous  : std_ulogic := 'X';
     variable LEVEL6_previous  : std_ulogic := 'X';
     variable LEVEL7_previous  : std_ulogic := 'X';

     -- Special variables to control flags
     variable hold_empty_low   : integer := 0;
     variable hold_eqth_high   : integer := 0;
     variable hold_geqth_high  : integer := 0;
     variable hold_full_low    : integer := 0;
     variable hold_empty_high  : integer := 0;
     variable hold_eqth_low    : integer := 0;
     variable hold_geqth_low   : integer := 0;
     variable WCLKS_re         : Time;
     variable WCLKS_fe         : Time;
     variable WCLKS_fe_prev    : Time;
     variable WB_re            : Time;
     variable RESET_re         : Time;


 begin -- process VITALBehavior

 if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

      VitalPeriodPulseCheck ( Pviol_RDB,
                              PeriodData_RDB,
                              RDB_ipd, "RDB",
                              0.0 ns,
                              tperiod_RDB,
                              tpw_RDB_posedge,
                              tpw_RDB_negedge,
                              (TO_X01(RBLKB) = '0') AND (TO_X01(RESET ) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9SA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RBLKB,
                              PeriodData_RBLKB,
                              RBLKB_ipd, "RBLKB",
                              0.0 ns,
                              tperiod_RBLKB,
                              tpw_RBLKB_posedge,
                              tpw_RBLKB_negedge,
                              (TO_X01(RDB) = '0') AND (TO_X01(RESET ) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9SA",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RESET,
                              PeriodData_RESET,
                              RESET_ipd, "RESET",
                              0.0 ns,
                              tpw_RESET_negedge,
                              0.0 ns,
                              tpw_RESET_negedge,
                              True,
                              InstancePath & "/FIFO256x9SA",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       -- recovery / removal check for WCLKS to RESET signal ;
       VitalRecoveryRemovalCheck ( Tviol_RESET_WCLKS_posedge,
                             Tmkr_RESET_WCLKS_posedge,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns,
                             trecovery_RESET_WCLKS_posedge_negedge,
                             thold_RESET_WCLKS_posedge_posedge,
                             TRUE,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'), 
                             '/',
                             InstancePath & "/FIFO256x9SA",
                             TRUE,
                             TRUE,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_posedge_posedge,
                             tsetup_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_posedge_posedge,
                             tsetup_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_posedge_posedge,
                             tsetup_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_posedge_posedge,
                             tsetup_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_posedge_posedge,
                             tsetup_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_posedge_posedge,
                             tsetup_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_posedge_posedge,
                             tsetup_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_posedge_posedge,
                             tsetup_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_posedge_posedge,
                             tsetup_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SA",
                             True,
                             True,
                             WARNING
                             );

   -- setup hold WEN, WBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_posedge_posedge,
                             tsetup_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SA",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_PARODD_WCLKS_posedge,
                             TmDt_PARODD_WCLKS_posedge,
                             PARODD_ipd, "PARODD",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_PARODD_WCLKS_posedge_posedge,
                             tsetup_PARODD_WCLKS_negedge_posedge,
                             thold_PARODD_WCLKS_posedge_posedge,
                             thold_PARODD_WCLKS_negedge_posedge,
                             ((TO_X01(RBint) = '0') AND (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/FIFO256x9SA",
                             True,
                             True,
                             WARNING
                             );

  --   Period of WCLK
      VitalPeriodPulseCheck ( Pviol_WCLKS,
                              PeriodData_WCLKS,
                              WCLKS_ipd, "WCLKS",
                              0.0 ns,
                              tperiod_WCLKS,
                              tpw_WCLKS_posedge,
                              tpw_WCLKS_negedge,
                              (TO_X01(WRB) = '0') AND (TO_X01(WBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9SA",
                              True,
                              True,
                              WARNING
                              );
 end if;

   ------------------------------------------------------------
   --               FIFO RESET                               --
   ------------------------------------------------------------

   if ( RESET_ipd'event and RESET_ipd = '0' ) then
       WADDR      := 0;
       RADDR      := 0;
       WADDR_wrap := 0;
       RADDR_wrap := 0;
       FULL_tmp   := '0';
       EMPTY_tmp  := '1';
       EQTH_tmp   := '0';
       GEQTH_tmp  := '0';
       WRITE_AT_PREV_EDGE <='0';
       --WPE_zd     := 'X';
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
       hold_full_low   := 0;
       hold_empty_high := 0;
       hold_eqth_low   := 0;
       hold_geqth_low  := 0;
   end if;

   if ( WCLKS_ipd'event and WCLKS_ipd = '1' ) then
     WCLKS_re := now;
   end if;
      
   if ( WBint'event and WBint = '1' ) then
     WB_re := now;
   end if;
      
   if ( RESET_ipd'event and RESET_ipd = '1' ) then
     RESET_re := now;
     if ( TO_X01 ( WCLKS_ipd ) = '1' ) then
       if ( WCLKS_re = WB_re ) then
         hold_full_low   := 1; -- until next reset
         hold_empty_high := 1;
         hold_eqth_low   := 1;
         hold_geqth_low  := 1;
       elsif ( TO_X01 ( WBint ) = '0' ) then
         EMPTY_zd        := '0';
         EQTH_zd         := '1';
         GEQTH_zd        := '1';
         hold_empty_low  := 1; -- until next WCLKS falling edge
         hold_eqth_high  := 1;
         hold_geqth_high := 1;
       elsif ( WCLKS_re < WB_re ) then
         EMPTY_zd        := '0';
         EQTH_zd         := '1';
         GEQTH_zd        := '1';
         hold_empty_low  := 1; -- until next WCLKS falling edge
         hold_eqth_high  := 1;
         hold_geqth_high := 1;
       elsif ( WB_re < WCLKS_re ) then
         hold_empty_low  := 0; -- expected behavior
         hold_eqth_high  := 0;
         hold_geqth_high := 0;
         hold_full_low   := 0;
         hold_empty_high := 0;
         hold_eqth_low   := 0;
         hold_geqth_low  := 0;
       end if;
     else
       hold_empty_low  := 0; -- expected behavior
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
       hold_full_low   := 0;
       hold_empty_high := 0;
       hold_eqth_low   := 0;
       hold_geqth_low  := 0;
     end if;
   end if;

   if ( WCLKS_ipd'event and WCLKS_ipd = '0' ) then
     WCLKS_fe_prev := WCLKS_fe;
     WCLKS_fe := now;
     if (( TO_X01 ( RESET_ipd ) = '1' ) and ( WCLKS_fe_prev < RESET_re )) then
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
     end if;
   end if;

   ------------------------------------------------------------
   -- WPE output                                              -
   ------------------------------------------------------------

   if ( PARODD_ipd'EVENT ) then
     RPE_zd := not RPE_zd;
     WPE_zd := not WPE_zd;
   end if;

   ------------------------------------------------------------
   --         WPE generating block                            -
   ------------------------------------------------------------

    if ( WCLKS_ipd'EVENT AND WCLKS_ipd = '1' ) then
      tmp_par := DI7_delayed XOR DI6_delayed XOR DI5_delayed XOR DI4_delayed XOR DI3_delayed XOR DI2_delayed XOR DI1_delayed XOR DI0_delayed;
      par_f    <= tmp_par ;
      tmp_par2 := ( tmp_par xor DI8_delayed );
      par_f2   <= tmp_par2;

      if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
          ( TO_X01 ( DI8_ipd )    = 'X' ) or
          ( TO_X01 ( DI7_ipd )    = 'X' ) or
          ( TO_X01 ( DI6_ipd )    = 'X' ) or
          ( TO_X01 ( DI5_ipd )    = 'X' ) or
          ( TO_X01 ( DI4_ipd )    = 'X' ) or
          ( TO_X01 ( DI3_ipd )    = 'X' ) or
          ( TO_X01 ( DI2_ipd )    = 'X' ) or
          ( TO_X01 ( DI1_ipd )    = 'X' ) or
          ( TO_X01 ( DI0_ipd )    = 'X' )
         ) then
        wpe_var  :=  'X';
      else
        if ( tmp_par2 /= PARODD_ipd ) then
          wpe_var  :=  '1';
        else
          wpe_var  :=  '0';
        end if;
      end if;
      RAM_di_int(8) := DI8_ipd;
      WPE_zd := wpe_var;
    end if;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

   if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
   end if; 

   -----------------------------------------------------------
   --    calculate the depth and levels                     --
   -----------------------------------------------------------

    temp :=((INT(LGDEP2_delayed)*4) + (INT(LGDEP1_delayed)*2) + 
           (INT(LGDEP0_delayed)*1));

    case temp is 
         when 0 => depth := 2;
         when 1 => depth := 4;
         when 2 => depth := 8;
         when 3 => depth := 16;
         when 4 => depth := 32;
         when 5 => depth := 64;
         when 6 => depth := 128;
         when 7 => depth := 256;
         when others => depth := 0;
    end case;

    -- thresh value

    thresh := (INT(LEVEL7_delayed)*128) + (INT(LEVEL6_delayed)*64) + 
               (INT(LEVEL5_delayed)*32) + (INT(LEVEL4_delayed)*16) + 
               (INT(LEVEL3_delayed)*8) + (INT(LEVEL2_delayed)*4) + 
               (INT(LEVEL1_delayed)*2) + (INT(LEVEL0_delayed)*1); 

    if ( thresh = 0 or thresh = 255 ) then
      assert false
        report " Illegal level configuration, LEVEL cannot be 0 or 255 "
        severity failure;
    end if;

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

   if ( TO_X01 ( WCLKS_ipd )='X' ) then
     if(RESET_delayed = '1') then
       if (WBint_delayed = '0') then
         if (TO_X01(WCLKS_previous) /= 'X') then
           assert false
           report ": WCLK unknown"
           severity Error;
         end if;
       end if;
     end if;
   elsif ( WCLKS_ipd'EVENT AND WCLKS_ipd = '1') AND (TO_X01(RESET_ipd) = '1') then
     WRITE_AT_PREV_EDGE <='0';
     case ( TO_X01 ( WBint_delayed )) is 
       when '1' =>
                null;
       when '0' => 
         if ( FULL_zd = '0' ) then 
           RAM_di_int ( 7 downto 0 ) := DI7_delayed & DI6_delayed & DI5_delayed & 
                                      DI4_delayed & DI3_delayed & DI2_delayed & 
                                      DI1_delayed & DI0_delayed;
           memory_array ( WADDR ) := RAM_di_int;
           WRITE_AT_PREV_EDGE <= '1';
           if ( WADDR < depth - 1 ) then
             WADDR := WADDR + 1;
           elsif ( WADDR  = depth - 1 ) then
             WADDR := 0;
             WADDR_wrap := 1 - WADDR_wrap;
           end if;
         end if;
       when others => 
         if ( TO_X01 ( WBint_previous ) /= 'X' ) then
           assert false
           report ": WBLKB or WRB unknown"
           severity Error;
         end if;
       end case;
     elsif (( WCLKS_ipd'EVENT AND WCLKS_ipd = '0' ) AND 
            ( TO_X01 ( RESET_delayed ) = '1'      )  AND 
            ( TO_X01 ( WRITE_AT_PREV_EDGE ) = '1' )
           ) then
        WRITE_AT_PREV_EDGE <='0';
        if ( WADDR = RADDR ) then
          if ( RADDR_wrap /= WADDR_wrap ) then
            FULL_tmp := '1';
            EMPTY_tmp :='0';
          end if;
        end if;
        if ( WADDR /= RADDR ) then
          EMPTY_tmp := '0';
        end if;
        if ( RADDR_wrap = WADDR_wrap ) then
          if ( WADDR - RADDR = thresh ) then
            EQTH_tmp := '1';
          else 
            EQTH_tmp := '0';
          end if;
          if ( WADDR - RADDR >= thresh ) then
            GEQTH_tmp := '1';
          else 
            GEQTH_tmp := '0';
          end if;
        else 
          if (( depth - RADDR + WADDR ) = thresh ) then
            EQTH_tmp := '1';
          else 
            EQTH_tmp := '0';
          end if;
          if (( depth - RADDR + WADDR ) >= thresh ) then
            GEQTH_tmp := '1';
          else 
            GEQTH_tmp := '0';
          end if;
        end if; 
      else
       null;
    end if;


  --------------------------------------------------------------------
  --          FIFO READ SECTION........                             --
  --------------------------------------------------------------------

  if ( TO_X01 ( RBint ) = 'X' ) then 
    if ( TO_X01 ( RESET_ipd ) /= '0' ) then 
      if ( TO_X01 ( RBint_previous ) /= 'X' ) then
        assert false
        report ": RDB or RBLKB unknown"
        severity error;
      end if;
     end if;
  elsif (( RBint'event AND TO_X01 ( RBint ) = '0' ) AND
         ( TO_X01 ( RESET_ipd ) /= '0'            )
        ) then
     if ( EMPTY_zd /= '1' ) then
       DO0_zd  := memory_array(RADDR)(0);
       DO1_zd  := memory_array(RADDR)(1);
       DO2_zd  := memory_array(RADDR)(2);
       DO3_zd  := memory_array(RADDR)(3);
       DO4_zd  := memory_array(RADDR)(4);
       DO5_zd  := memory_array(RADDR)(5);
       DO6_zd  := memory_array(RADDR)(6);
       DO7_zd  := memory_array(RADDR)(7);
       DO8_zd  := memory_array(RADDR)(8);
     if ( RADDR < depth - 1 ) then
       RADDR := RADDR + 1;
     else
       RADDR :=(RADDR +1) mod  depth;
       RADDR_wrap :=1 - RADDR_wrap;
     end if;
             do_par  :=DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR
                       DO3_zd XOR DO2_zd XOR DO1_zd XOR DO0_zd;
             par_f <= do_par;
             if (do_par = 'X') then
               RPE_zd := 'X';
             elsif (do_par /= PARODD_ipd) then
               RPE_zd := '1';
             else
               RPE_zd :=  '0';
             end if;
     end if;
  else 
   null;
  end if;
  if (( RBint'event and TO_X01 ( RBint ) ='1') AND 
      ( TO_X01 ( RESET_ipd ) /= '0'          ) AND
      ( EMPTY_zd /= '1'                      )
     ) then
    if ( RADDR = WADDR ) then
      if ( RADDR_wrap = WADDR_wrap ) then
        EMPTY_tmp := '1';
        FULL_tmp   :=  '0';
      end if;
    end if;
    if ( RADDR /= WADDR ) then
      FULL_tmp  := '0';
    end if;
    if ( WADDR_wrap = RADDR_wrap ) then
      if (( WADDR - RADDR ) = thresh ) then
        EQTH_tmp := '1';
      else
        EQTH_tmp := '0';
      end if;
      if (( WADDR - RADDR ) >= thresh ) then
        GEQTH_tmp := '1';
      else
        GEQTH_tmp := '0';
      end if;
    else 
      if (( depth + WADDR - RADDR ) = thresh ) then
        EQTH_tmp := '1';
      else
        EQTH_tmp := '0';
      end if;
      if (( depth + WADDR - RADDR ) >= thresh ) then
        GEQTH_tmp := '1';
      else
        GEQTH_tmp := '0';
      end if;
    end if;
  end if;

   -- Mimic odd silicon flag behavior coming out of RESET with WB low
   
   if ( hold_full_low = 1 ) then
     FULL_zd := '0';
   else
     FULL_zd := FULL_tmp;
   end if;

   if ( hold_empty_low = 1 ) then
     EMPTY_zd := '0';
   elsif ( hold_empty_high = 1 ) then
     EMPTY_zd := '1';
   else
     EMPTY_zd := EMPTY_tmp;
   end if;

   if ( hold_eqth_high = 1 ) then
     EQTH_zd := '1';
   elsif ( hold_eqth_low = 1 ) then
     EQTH_zd := '0';
   else
     EQTH_zd := EQTH_tmp;
   end if;

   -- If LEVEL greater than DEPTH then GEQTH mimics FULL
   
   if ( hold_geqth_high = 1 ) then
     GEQTH_zd := '1';
   elsif ( hold_geqth_low = 1 ) then
     GEQTH_zd := '0';
   else
     if ( thresh > depth ) then
       GEQTH_zd := FULL_zd;
     else
       GEQTH_zd := GEQTH_tmp;
     end if;
   end if;

  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       WCLKS_previous  := WCLKS_ipd;
       RBint_previous   := RBint;
       WBint_previous   := WBint_delayed;
       WBint_delayed    := WBint;
       DI0_delayed      := DI0_ipd;
       DI1_delayed      := DI1_ipd;
       DI2_delayed      := DI2_ipd;
       DI3_delayed      := DI3_ipd;
       DI4_delayed      := DI4_ipd;
       DI5_delayed      := DI5_ipd;
       DI6_delayed      := DI6_ipd;
       DI7_delayed      := DI7_ipd;
       DI8_delayed      := DI8_ipd;
       LGDEP0_previous  := LGDEP0_delayed;
       LGDEP0_delayed   := LGDEP0_ipd;
       LGDEP1_previous  := LGDEP1_delayed;
       LGDEP1_delayed   := LGDEP1_ipd;
       LGDEP2_previous  := LGDEP2_delayed;
       LGDEP2_delayed   := LGDEP2_ipd;
       LEVEL0_previous  := LEVEL0_delayed;
       LEVEL0_delayed   := LEVEL0_ipd;
       LEVEL1_previous  := LEVEL1_delayed;
       LEVEL1_delayed   := LEVEL1_ipd;
       LEVEL2_previous  := LEVEL2_delayed;
       LEVEL2_delayed   := LEVEL2_ipd;
       LEVEL3_previous  := LEVEL3_delayed;
       LEVEL3_delayed   := LEVEL3_ipd;
       LEVEL4_previous  := LEVEL4_delayed;
       LEVEL4_delayed   := LEVEL4_ipd;
       LEVEL5_previous  := LEVEL5_delayed;
       LEVEL5_delayed   := LEVEL5_ipd;
       LEVEL6_previous  := LEVEL6_delayed;
       LEVEL6_delayed   := LEVEL6_ipd;
       LEVEL7_previous  := LEVEL7_delayed;
       LEVEL7_delayed   := LEVEL7_ipd;
       PARODD_previous  := PARODD_delayed; 
       PARODD_delayed   := PARODD_ipd;
       RESET_previous   := RESET_delayed; 
       RESET_delayed    := RESET_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
             OutSignal     => DOS,
             GlitchData    => DOS_GlitchData,
             OutSignalName => "DOS",
             OutTemp       => DOS_zd,

             Paths =>   (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
           OutSignal     => WPE,
           GlitchData    => WPE_GlitchData,
           OutSignalName => "WPE",
           OutTemp       => WPE_zd,
           Paths =>   (0  => (WCLKS_ipd'last_event,
                             VitalExtendToFillDelay(tpd_WCLKS_WPE), true),
                       1 => (PARODD_ipd'last_event,
                             VitalExtendToFillDelay(tpd_PARODD_WPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO0), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO0), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO1), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO1), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO2), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO2), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO3), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO3), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO4), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO4), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO5), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO5), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO6), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO6), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO7), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO7), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO8), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO8), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => RPE,
           GlitchData    => RPE_GlitchData,
           OutSignalName => "RPE",
           OutTemp       => RPE_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_RPE), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_RPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => FULL,
           GlitchData    => FULL_GlitchData,
           OutSignalName => "FULL",
           OutTemp       => FULL_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_FULL), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_FULL), true),
                       2 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_FULL), true),
                       3 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_FULL), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EMPTY,
           GlitchData    => EMPTY_GlitchData,
           OutSignalName => "EMPTY",
           OutTemp       => EMPTY_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EMPTY), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_EMPTY), true),
                       2 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_EMPTY), true),
                       3 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_EMPTY), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EQTH,
           GlitchData    => EQTH_GlitchData,
           OutSignalName => "EQTH",
           OutTemp       => EQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EQTH), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_EQTH), true),
                       2 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_EQTH), true),
                       3 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_EQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => GEQTH,
           GlitchData    => GEQTH_GlitchData,
           OutSignalName => "GEQTH",
           OutTemp       => GEQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_GEQTH), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_GEQTH), true),
                       2 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_GEQTH), true),
                       3 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_GEQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );


   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

LIBRARY a500k;
USE a500k.all;

entity FIFO256x9SAP is 
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_RBLKB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RBLKB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RDB_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tpw_RDB_posedge         : VitalDelayType        := 0.000 ns;
 	tpw_RDB_negedge         : VitalDelayType        := 0.000 ns;
 	tperiod_RDB             : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_posedge       : VitalDelayType        := 0.000 ns;
 	tpw_RBLKB_negedge       : VitalDelayType        := 0.000 ns;
 	tperiod_RBLKB           : VitalDelayType        := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_WCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_WCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;

        -- WCLK falling edge setup to RESET rising edge 
 	trecovery_RESET_WCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_WCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- WCLK rising  edge hold to RESET rising edge 
	thold_RESET_WCLKS_posedge_posedge             : VitalDelayType := 0.00 ns;
	thold_RESET_WCLKS_posedge_negedge             : VitalDelayType := 0.00 ns;
	tpw_WCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        WCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');


ATTRIBUTE VITAL_LEVEL0 OF FIFO256x9SAP : entity IS True ;
END FIFO256x9SAP;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of FIFO256x9SAP is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal LGDEP0_ipd : std_ulogic := 'X';
   signal LGDEP1_ipd : std_ulogic := 'X';
   signal LGDEP2_ipd : std_ulogic := 'X';
   signal LEVEL0_ipd : std_ulogic := 'X';
   signal LEVEL1_ipd : std_ulogic := 'X';
   signal LEVEL2_ipd : std_ulogic := 'X';
   signal LEVEL3_ipd : std_ulogic := 'X';
   signal LEVEL4_ipd : std_ulogic := 'X';
   signal LEVEL5_ipd : std_ulogic := 'X';
   signal LEVEL6_ipd : std_ulogic := 'X';
   signal LEVEL7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal RESET_ipd  : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal WCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

   -- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic := 'X';
   signal par_f2     : std_logic := 'X';

   signal WRITE_AT_PREV_EDGE : std_logic := '0';
   signal READ_AT_PREV_EDGE  : std_logic := '0';

   begin  --  VITAL_ACT

   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (LGDEP0_ipd, LGDEP0, VitalExtendToFillDelay(tipd_LGDEP0));
   VitalWireDelay (LGDEP1_ipd, LGDEP1, VitalExtendToFillDelay(tipd_LGDEP1));
   VitalWireDelay (LGDEP2_ipd, LGDEP2, VitalExtendToFillDelay(tipd_LGDEP2));
   VitalWireDelay (LEVEL0_ipd, LEVEL0, VitalExtendToFillDelay(tipd_LEVEL0));
   VitalWireDelay (LEVEL1_ipd, LEVEL1, VitalExtendToFillDelay(tipd_LEVEL1));
   VitalWireDelay (LEVEL2_ipd, LEVEL2, VitalExtendToFillDelay(tipd_LEVEL2));
   VitalWireDelay (LEVEL3_ipd, LEVEL3, VitalExtendToFillDelay(tipd_LEVEL3));
   VitalWireDelay (LEVEL4_ipd, LEVEL4, VitalExtendToFillDelay(tipd_LEVEL4));
   VitalWireDelay (LEVEL5_ipd, LEVEL5, VitalExtendToFillDelay(tipd_LEVEL5));
   VitalWireDelay (LEVEL6_ipd, LEVEL6, VitalExtendToFillDelay(tipd_LEVEL6));
   VitalWireDelay (LEVEL7_ipd, LEVEL7, VitalExtendToFillDelay(tipd_LEVEL7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RESET_ipd, RESET, VitalExtendToFillDelay(tipd_RESET));
   VitalWireDelay (WCLKS_ipd, WCLKS, VitalExtendToFillDelay(tipd_WCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

   ---------------------------------------------------------------
   --                  Behavior Section                         --
   ---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);

    VITALBehavior : process (
                          LEVEL0_ipd, LEVEL1_ipd, LEVEL2_ipd, LEVEL3_ipd, LEVEL4_ipd, LEVEL5_ipd, LEVEL6_ipd, LEVEL7_ipd, 
                          LGDEP0_ipd, LGDEP1_ipd, LGDEP2_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          WCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd, RESET_ipd
                          )

     -- some internal veriable declaration
     variable RAM_di_int   : std_logic_vector(8 downto 0);
     variable memory_array : MEM_TYPE  := (others =>(others => 'X'));
     variable do_par       : std_logic := 'X';
     variable tmp_par      : std_logic := 'X';
     variable tmp_par2     : std_logic := 'X';
     variable wpe_var      : std_logic := 'X';
     variable temp         : integer   := 0;
     variable thresh       : integer   := 0;
     variable depth        : integer   := 0;
     variable WADDR        : integer   := 0;
     variable WADDR_wrap   : integer   := 0;
     variable RADDR        : integer   := 0;
     variable RADDR_wrap   : integer   := 0;

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     --  Read Timing Check Results
     variable PeriodData_RESET           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET                : X01                 := '0';
     variable PeriodData_RDB             : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RDB                  : X01                 := '0';
     variable PeriodData_RBLKB           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RBLKB                : X01                 := '0';
     variable Tviol_DI0_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI0_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI1_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI2_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI3_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI4_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI5_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI6_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI7_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI8_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_PARODD_WCLKS_posedge : X01                 := '0';
     variable TmDt_PARODD_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_WCLKS_posedge    : X01                 := '0';
     variable TmDt_WRB_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_WCLKS_posedge  : X01                 := '0';
     variable TmDt_WBLKB_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_WCLKS_posedge  : X01                 := '0';
     variable Tmkr_RESET_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WCLKS                : X01                 := '0';

     -- functional Results


     variable DO0_zd   : std_ulogic;
     variable DO1_zd   : std_ulogic;
     variable DO2_zd   : std_ulogic;
     variable DO3_zd   : std_ulogic;
     variable DO4_zd   : std_ulogic;
     variable DO5_zd   : std_ulogic;
     variable DO6_zd   : std_ulogic;
     variable DO7_zd   : std_ulogic;
     variable DO8_zd   : std_ulogic;
     variable RPE_zd   : std_ulogic;
     variable WPE_zd   : std_ulogic;
     variable DOS_zd   : std_ulogic;
     variable FULL_zd  : std_ulogic;
     variable EMPTY_zd : std_ulogic;
     variable EQTH_zd  : std_ulogic;
     variable GEQTH_zd : std_ulogic;
     variable FULL_tmp  : std_ulogic;
     variable EMPTY_tmp : std_ulogic;
     variable EQTH_tmp  : std_ulogic;
     variable GEQTH_tmp : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData   : VitalGlitchDataType;
     variable DO1_GlitchData   : VitalGlitchDataType;
     variable DO2_GlitchData   : VitalGlitchDataType;
     variable DO3_GlitchData   : VitalGlitchDataType;
     variable DO4_GlitchData   : VitalGlitchDataType;
     variable DO5_GlitchData   : VitalGlitchDataType;
     variable DO6_GlitchData   : VitalGlitchDataType;
     variable DO7_GlitchData   : VitalGlitchDataType;
     variable DO8_GlitchData   : VitalGlitchDataType;
     variable DOS_GlitchData   : VitalGlitchDataType;
     variable FULL_GlitchData  : VitalGlitchDataType;
     variable EMPTY_GlitchData : VitalGlitchDataType;
     variable EQTH_GlitchData  : VitalGlitchDataType;
     variable GEQTH_GlitchData : VitalGlitchDataType;

     -- last value variables
     variable WCLKS_previous   : std_ulogic := 'X';
     variable RBint_previous   : std_ulogic := 'X';
     variable WBint_delayed    : std_ulogic := 'X';
     variable WBint_previous   : std_ulogic := 'X';
     variable DIS_previous     : std_ulogic := 'X';
     variable RESET_previous   : std_ulogic := 'X';
     variable RESET_delayed    : std_ulogic := 'X';
     variable PARODD_previous  : std_ulogic := 'X';
     variable PARODD_delayed   : std_ulogic := 'X';
     variable DI0_delayed      : std_ulogic := 'X';
     variable DI1_delayed      : std_ulogic := 'X';
     variable DI2_delayed      : std_ulogic := 'X';
     variable DI3_delayed      : std_ulogic := 'X';
     variable DI4_delayed      : std_ulogic := 'X';
     variable DI5_delayed      : std_ulogic := 'X';
     variable DI6_delayed      : std_ulogic := 'X';
     variable DI7_delayed      : std_ulogic := 'X';
     variable DI8_delayed      : std_ulogic := 'X';
     variable DI0_previous     : std_ulogic := 'X';
     variable DI1_previous     : std_ulogic := 'X';
     variable DI2_previous     : std_ulogic := 'X';
     variable DI3_previous     : std_ulogic := 'X';
     variable DI4_previous     : std_ulogic := 'X';
     variable DI5_previous     : std_ulogic := 'X';
     variable DI6_previous     : std_ulogic := 'X';
     variable DI7_previous     : std_ulogic := 'X';
     variable DI8_previous     : std_ulogic := 'X';
     variable LGDEP0_delayed   : std_ulogic := 'X';
     variable LGDEP1_delayed   : std_ulogic := 'X';
     variable LGDEP2_delayed   : std_ulogic := 'X';
     variable LGDEP0_previous  : std_ulogic := 'X';
     variable LGDEP1_previous  : std_ulogic := 'X';
     variable LGDEP2_previous  : std_ulogic := 'X';
     variable LEVEL0_delayed   : std_ulogic := 'X';
     variable LEVEL1_delayed   : std_ulogic := 'X';
     variable LEVEL2_delayed   : std_ulogic := 'X';
     variable LEVEL3_delayed   : std_ulogic := 'X';
     variable LEVEL4_delayed   : std_ulogic := 'X';
     variable LEVEL5_delayed   : std_ulogic := 'X';
     variable LEVEL6_delayed   : std_ulogic := 'X';
     variable LEVEL7_delayed   : std_ulogic := 'X';
     variable LEVEL0_previous  : std_ulogic := 'X';
     variable LEVEL1_previous  : std_ulogic := 'X';
     variable LEVEL2_previous  : std_ulogic := 'X';
     variable LEVEL3_previous  : std_ulogic := 'X';
     variable LEVEL4_previous  : std_ulogic := 'X';
     variable LEVEL5_previous  : std_ulogic := 'X';
     variable LEVEL6_previous  : std_ulogic := 'X';
     variable LEVEL7_previous  : std_ulogic := 'X';

     -- Special variables to control flags
     variable hold_empty_low   : integer := 0;
     variable hold_eqth_high   : integer := 0;
     variable hold_geqth_high  : integer := 0;
     variable hold_full_low    : integer := 0;
     variable hold_empty_high  : integer := 0;
     variable hold_eqth_low    : integer := 0;
     variable hold_geqth_low   : integer := 0;

     variable WCLKS_re         : Time;
     variable WCLKS_fe         : Time;
     variable WCLKS_fe_prev    : Time;
     variable WB_re            : Time;
     variable RESET_re         : Time;

 begin -- process VITALBehavior

 if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

      VitalPeriodPulseCheck ( Pviol_RDB,
                              PeriodData_RDB,
                              RDB_ipd, "RDB",
                              0.0 ns,
                              tperiod_RDB,
                              tpw_RDB_posedge,
                              tpw_RDB_negedge,
                              (TO_X01(RBLKB) = '0') AND (TO_X01(RESET ) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9SAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RBLKB,
                              PeriodData_RBLKB,
                              RBLKB_ipd, "RBLKB",
                              0.0 ns,
                              tperiod_RBLKB,
                              tpw_RBLKB_posedge,
                              tpw_RBLKB_negedge,
                              (TO_X01(RDB) = '0') AND (TO_X01(RESET ) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9SAP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RESET,
                              PeriodData_RESET,
                              RESET_ipd, "RESET",
                              0.0 ns,
                              tpw_RESET_negedge,
                              0.0 ns,
                              tpw_RESET_negedge,
                              True,
                              InstancePath & "/FIFO256x9SAP",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       -- recovery / removal check for WCLKS to RESET signal ;
       VitalRecoveryRemovalCheck ( Tviol_RESET_WCLKS_posedge,
                             Tmkr_RESET_WCLKS_posedge,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns,
                             trecovery_RESET_WCLKS_posedge_negedge,
                             thold_RESET_WCLKS_posedge_posedge,
                             TRUE,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'), 
                             '/',
                             InstancePath & "/FIFO256x9SAP",
                             TRUE,
                             TRUE,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_posedge_posedge,
                             tsetup_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_posedge_posedge,
                             tsetup_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_posedge_posedge,
                             tsetup_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_posedge_posedge,
                             tsetup_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_posedge_posedge,
                             tsetup_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_posedge_posedge,
                             tsetup_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_posedge_posedge,
                             tsetup_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_posedge_posedge,
                             tsetup_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_posedge_posedge,
                             tsetup_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SAP",
                             True,
                             True,
                             WARNING
                             );

   -- setup hold WEN, WBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_posedge_posedge,
                             tsetup_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SAP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_PARODD_WCLKS_posedge,
                             TmDt_PARODD_WCLKS_posedge,
                             PARODD_ipd, "PARODD",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_PARODD_WCLKS_posedge_posedge,
                             tsetup_PARODD_WCLKS_negedge_posedge,
                             thold_PARODD_WCLKS_posedge_posedge,
                             thold_PARODD_WCLKS_negedge_posedge,
                             ((TO_X01(RBint) = '0') AND (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/FIFO256x9SAP",
                             True,
                             True,
                             WARNING
                             );

  --   Period of WCLK
      VitalPeriodPulseCheck ( Pviol_WCLKS,
                              PeriodData_WCLKS,
                              WCLKS_ipd, "WCLKS",
                              0.0 ns,
                              tperiod_WCLKS,
                              tpw_WCLKS_posedge,
                              tpw_WCLKS_negedge,
                              (TO_X01(WRB) = '0') AND (TO_X01(WBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9SAP",
                              True,
                              True,
                              WARNING
                              );
 end if;

   ------------------------------------------------------------
   --               FIFO RESET                               --
   ------------------------------------------------------------

   if ( RESET_ipd'event and RESET_ipd = '0' ) then
       WADDR      := 0;
       RADDR      := 0;
       WADDR_wrap := 0;
       RADDR_wrap := 0;
       FULL_tmp   := '0';
       EMPTY_tmp  := '1';
       EQTH_tmp   := '0';
       GEQTH_tmp  := '0';
       WRITE_AT_PREV_EDGE <='0';
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
       hold_full_low   := 0;
       hold_empty_high := 0;
       hold_eqth_low   := 0;
       hold_geqth_low  := 0;
   end if;

   if ( WCLKS_ipd'event and WCLKS_ipd = '1' ) then
     WCLKS_re := now;
   end if;
      
   if ( WBint'event and WBint = '1' ) then
     WB_re := now;
   end if;
      
   if ( RESET_ipd'event and RESET_ipd = '1' ) then
     RESET_re := now;
     if ( TO_X01 ( WCLKS_ipd ) = '1' ) then
       if ( WCLKS_re = WB_re ) then
         hold_full_low   := 1; -- until next reset
         hold_empty_high := 1;
         hold_eqth_low   := 1;
         hold_geqth_low  := 1;
       elsif ( TO_X01 ( WBint ) = '0' ) then
         EMPTY_zd        := '0';
         EQTH_zd         := '1';
         GEQTH_zd        := '1';
         hold_empty_low  := 1; -- until next WCLKS falling edge
         hold_eqth_high  := 1;
         hold_geqth_high := 1;
       elsif ( WCLKS_re < WB_re ) then
         EMPTY_zd        := '0';
         EQTH_zd         := '1';
         GEQTH_zd        := '1';
         hold_empty_low  := 1; -- until next WCLKS falling edge
         hold_eqth_high  := 1;
         hold_geqth_high := 1;
       elsif ( WB_re < WCLKS_re ) then
         hold_empty_low  := 0; -- expected behavior
         hold_eqth_high  := 0;
         hold_geqth_high := 0;
         hold_full_low   := 0;
         hold_empty_high := 0;
         hold_eqth_low   := 0;
         hold_geqth_low  := 0;
       end if;
     else
       hold_empty_low  := 0; -- expected behavior
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
       hold_full_low   := 0;
       hold_empty_high := 0;
       hold_eqth_low   := 0;
       hold_geqth_low  := 0;
     end if;
   end if;

   if ( WCLKS_ipd'event and WCLKS_ipd = '0' ) then
     WCLKS_fe_prev := WCLKS_fe;
     WCLKS_fe := now;
     if (( TO_X01 ( RESET_ipd ) = '1' ) and ( WCLKS_fe_prev < RESET_re )) then
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
     end if;
   end if;


   ------------------------------------------------------------
   --         WPE generating block                            -
   ------------------------------------------------------------

    if (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      tmp_par  := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;
      par_f  <= tmp_par ;
      if (tmp_par /= PARODD_ipd) then
        wpe_var  :=  '1';
      else
        wpe_var  :=  '0';
      end if;
      RAM_di_int(8) := wpe_var;
      WPE_zd := wpe_var;
    end if;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

   if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
   end if; 

   -----------------------------------------------------------
   --    calculate the depth and levels                     --
   -----------------------------------------------------------

    temp :=((INT(LGDEP2_delayed)*4) + (INT(LGDEP1_delayed)*2) + 
           (INT(LGDEP0_delayed)*1));

    case temp is 
         when 0 => depth := 2;
         when 1 => depth := 4;
         when 2 => depth := 8;
         when 3 => depth := 16;
         when 4 => depth := 32;
         when 5 => depth := 64;
         when 6 => depth := 128;
         when 7 => depth := 256;
         when others => depth := 0;
    end case;

    -- thresh value

    thresh := (INT(LEVEL7_delayed)*128) + (INT(LEVEL6_delayed)*64) + 
               (INT(LEVEL5_delayed)*32) + (INT(LEVEL4_delayed)*16) + 
               (INT(LEVEL3_delayed)*8) + (INT(LEVEL2_delayed)*4) + 
               (INT(LEVEL1_delayed)*2) + (INT(LEVEL0_delayed)*1); 

    if ( thresh = 0 or thresh = 255 ) then
      assert false
        report " Illegal level configuration, LEVEL cannot be 0 or 255 "
        severity failure;
    end if;

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

   if(TO_X01(WCLKS_ipd)='X') then
    if(RESET_delayed = '1') then
     if (WBint_delayed = '0') then
      if (TO_X01(WCLKS_previous) /= 'X') then
        assert false
        report ": WCLK unknown"
        severity Error;
      end if;
     end if;
    end if;
   elsif (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') AND (TO_X01(RESET_ipd) = '1')then
     WRITE_AT_PREV_EDGE <='0';
     case (TO_X01(WBint_delayed)) is 
      when '1' =>
                null;
      when '0' => 
         if(FULL_zd = '0') then 
         RAM_di_int(7 downto 0) := DI7_delayed & DI6_delayed & DI5_delayed & 
                                    DI4_delayed & DI3_delayed & DI2_delayed & 
                                    DI1_delayed & DI0_delayed;
         memory_array(WADDR) := RAM_di_int;
         WRITE_AT_PREV_EDGE <='1';
         if(WADDR <depth-1  ) then
           WADDR := WADDR + 1;
         elsif( WADDR  = depth-1) then
           WADDR := 0;
           WADDR_wrap := 1 - WADDR_wrap;
         end if;
        end if;
       when others => 
        if (TO_X01(WBint_previous) /= 'X') then
          assert false
          report ": WBLKB or WRB unknown"
          severity Error;
          end if;
        end case;
     elsif(WCLKS_ipd'EVENT AND WCLKS_ipd = '0')  AND (TO_X01(RESET_delayed) = '1') AND (TO_X01(WRITE_AT_PREV_EDGE) = '1')then
        WRITE_AT_PREV_EDGE <='0';
        if(WADDR   = RADDR ) then
         if(RADDR_wrap /= WADDR_wrap) then
          FULL_tmp := '1';
          EMPTY_tmp :='0';
         end if;
        end if;
        if(WADDR   /= RADDR ) then
          EMPTY_tmp := '0';
        end if;
          if(RADDR_wrap = WADDR_wrap) then
            if(WADDR - RADDR = thresh ) then
               EQTH_tmp := '1';
            else 
               EQTH_tmp := '0';
            end if;
            if(WADDR - RADDR >= thresh ) then
                GEQTH_tmp := '1';
            else 
                GEQTH_tmp := '0';
            end if;
          else 
           if((depth -RADDR + WADDR) = thresh ) then
               EQTH_tmp := '1';
            else 
               EQTH_tmp := '0';
            end if;
            if((depth -RADDR + WADDR) >= thresh ) then
                GEQTH_tmp := '1';
            else 
                GEQTH_tmp := '0';
            end if;
           end if; 
      else
       null;
    end if;


  --------------------------------------------------------------------
  --          FIFO READ SECTION........                             --
  --------------------------------------------------------------------

  if(TO_X01(RBint) = 'X') then 
    if(TO_X01(RESET_ipd) /= '0') then 
      if(TO_X01(RBint_previous) /= 'X') then
        assert false
        report ": RDB or RBLKB unknown"
        severity error;
      end if;
     end if;
  elsif (( RBint'event AND TO_X01 ( RBint ) = '0' ) AND
         ( TO_X01 ( RESET_ipd ) /= '0'            )
        ) then
     if(EMPTY_zd /= '1') then
           DO0_zd  := memory_array(RADDR)(0);
           DO1_zd  := memory_array(RADDR)(1);
           DO2_zd  := memory_array(RADDR)(2);
           DO3_zd  := memory_array(RADDR)(3);
           DO4_zd  := memory_array(RADDR)(4);
           DO5_zd  := memory_array(RADDR)(5);
           DO6_zd  := memory_array(RADDR)(6);
           DO7_zd  := memory_array(RADDR)(7);
           DO8_zd  := memory_array(RADDR)(8);
     if(RADDR <depth-1  ) then
        RADDR := RADDR + 1;
     else
        RADDR :=(RADDR +1) mod  depth;
        RADDR_wrap :=1 - RADDR_wrap;
     end if;
             do_par  :=DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR
                       DO3_zd XOR DO2_zd XOR DO1_zd XOR DO0_zd;
             par_f <= do_par;
             if (do_par = 'X') then
               RPE_zd := 'X';
             elsif (do_par /= PARODD_ipd) then
               RPE_zd := '1';
             else
               RPE_zd :=  '0';
             end if;
     end if;
  else 
   null;
  end if;
  if (( RBint'event and TO_X01 ( RBint ) ='1') AND 
      ( TO_X01 ( RESET_ipd ) /= '0'          ) AND
      ( EMPTY_zd /= '1'                      )
     ) then
    if(RADDR = WADDR ) then
     if(RADDR_wrap = WADDR_wrap) then
       EMPTY_tmp := '1';
       FULL_tmp   :=  '0';
     end if;
    end if;
    if(RADDR /= WADDR ) then
     FULL_tmp  := '0';
    end if;
     if(WADDR_wrap = RADDR_wrap ) then
      if((WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
      else
       EQTH_tmp := '0';
      end if;
      if((WADDR - RADDR) >= thresh ) then
       GEQTH_tmp := '1';
      else
       GEQTH_tmp := '0';
      end if;
    else 
     if((depth + WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((depth + WADDR - RADDR) >= thresh ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    end if;
   end if;


   -- Mimic odd silicon flag behavior coming out of RESET with WB low
   
   if ( hold_full_low = 1 ) then
     FULL_zd := '0';
   else
     FULL_zd := FULL_tmp;
   end if;

   if ( hold_empty_low = 1 ) then
     EMPTY_zd := '0';
   elsif ( hold_empty_high = 1 ) then
     EMPTY_zd := '1';
   else
     EMPTY_zd := EMPTY_tmp;
   end if;

   if ( hold_eqth_high = 1 ) then
     EQTH_zd := '1';
   elsif ( hold_eqth_low = 1 ) then
     EQTH_zd := '0';
   else
     EQTH_zd := EQTH_tmp;
   end if;

   -- If LEVEL greater than DEPTH then GEQTH mimics FULL
   
   if ( hold_geqth_high = 1 ) then
     GEQTH_zd := '1';
   elsif ( hold_geqth_low = 1 ) then
     GEQTH_zd := '0';
   else
     if ( thresh > depth ) then
       GEQTH_zd := FULL_zd;
     else
       GEQTH_zd := GEQTH_tmp;
     end if;
   end if;


  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       WCLKS_previous  := WCLKS_ipd;
       RBint_previous   := RBint;
       WBint_previous   := WBint_delayed;
       WBint_delayed    := WBint;
       DI0_delayed      := DI0_ipd;
       DI1_delayed      := DI1_ipd;
       DI2_delayed      := DI2_ipd;
       DI3_delayed      := DI3_ipd;
       DI4_delayed      := DI4_ipd;
       DI5_delayed      := DI5_ipd;
       DI6_delayed      := DI6_ipd;
       DI7_delayed      := DI7_ipd;
       DI8_delayed      := DI8_ipd;
       LGDEP0_previous  := LGDEP0_delayed;
       LGDEP0_delayed   := LGDEP0_ipd;
       LGDEP1_previous  := LGDEP1_delayed;
       LGDEP1_delayed   := LGDEP1_ipd;
       LGDEP2_previous  := LGDEP2_delayed;
       LGDEP2_delayed   := LGDEP2_ipd;
       LEVEL0_previous  := LEVEL0_delayed;
       LEVEL0_delayed   := LEVEL0_ipd;
       LEVEL1_previous  := LEVEL1_delayed;
       LEVEL1_delayed   := LEVEL1_ipd;
       LEVEL2_previous  := LEVEL2_delayed;
       LEVEL2_delayed   := LEVEL2_ipd;
       LEVEL3_previous  := LEVEL3_delayed;
       LEVEL3_delayed   := LEVEL3_ipd;
       LEVEL4_previous  := LEVEL4_delayed;
       LEVEL4_delayed   := LEVEL4_ipd;
       LEVEL5_previous  := LEVEL5_delayed;
       LEVEL5_delayed   := LEVEL5_ipd;
       LEVEL6_previous  := LEVEL6_delayed;
       LEVEL6_delayed   := LEVEL6_ipd;
       LEVEL7_previous  := LEVEL7_delayed;
       LEVEL7_delayed   := LEVEL7_ipd;
       PARODD_previous  := PARODD_delayed; 
       PARODD_delayed   := PARODD_ipd;
       RESET_previous   := RESET_delayed; 
       RESET_delayed    := RESET_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
             OutSignal     => DOS,
             GlitchData    => DOS_GlitchData,
             OutSignalName => "DOS",
             OutTemp       => DOS_zd,

             Paths =>   (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO0), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO0), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO1), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO1), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO2), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO2), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO3), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO3), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO4), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO4), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO5), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO5), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO6), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO6), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO7), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO7), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths =>   (0 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_DO8), true),
                       1 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_DO8), true),
                       2 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => FULL,
           GlitchData    => FULL_GlitchData,
           OutSignalName => "FULL",
           OutTemp       => FULL_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_FULL), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_FULL), true),
                       2 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_FULL), true),
                       3 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_FULL), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EMPTY,
           GlitchData    => EMPTY_GlitchData,
           OutSignalName => "EMPTY",
           OutTemp       => EMPTY_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EMPTY), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_EMPTY), true),
                       2 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_EMPTY), true),
                       3 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_EMPTY), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EQTH,
           GlitchData    => EQTH_GlitchData,
           OutSignalName => "EQTH",
           OutTemp       => EQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EQTH), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_EQTH), true),
                       2 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_EQTH), true),
                       3 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_EQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => GEQTH,
           GlitchData    => GEQTH_GlitchData,
           OutSignalName => "GEQTH",
           OutTemp       => GEQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_GEQTH), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_GEQTH), true),
                       2 => (RDB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RDB_GEQTH), true),
                       3 => (RBLKB_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RBLKB_GEQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );


   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

LIBRARY a500k;
USE a500k.all;

entity FIFO256x9SST is 
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_PARODD_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_WCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_WCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;

        -- WCLK falling edge setup to RESET rising edge 
 	trecovery_RESET_WCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_WCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- WCLK rising  edge hold to RESET rising edge 
	thold_RESET_WCLKS_posedge_posedge             : VitalDelayType := 0.00 ns;
	thold_RESET_WCLKS_posedge_negedge             : VitalDelayType := 0.00 ns;
	tpw_WCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        WPE    :  OUT STD_LOGIC := 'X';
        RPE    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        WCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');


ATTRIBUTE VITAL_LEVEL0 OF FIFO256x9SST : entity IS True ;
END FIFO256x9SST;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of FIFO256x9SST is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal LGDEP0_ipd : std_ulogic := 'X';
   signal LGDEP1_ipd : std_ulogic := 'X';
   signal LGDEP2_ipd : std_ulogic := 'X';
   signal LEVEL0_ipd : std_ulogic := 'X';
   signal LEVEL1_ipd : std_ulogic := 'X';
   signal LEVEL2_ipd : std_ulogic := 'X';
   signal LEVEL3_ipd : std_ulogic := 'X';
   signal LEVEL4_ipd : std_ulogic := 'X';
   signal LEVEL5_ipd : std_ulogic := 'X';
   signal LEVEL6_ipd : std_ulogic := 'X';
   signal LEVEL7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal RESET_ipd  : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal WCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

   -- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic := 'X';
   signal par_f2     : std_logic := 'X';

   signal WRITE_AT_PREV_EDGE : std_logic := '0';
   signal READ_AT_PREV_EDGE  : std_logic := '0';

   begin  --  VITAL_ACT

   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (LGDEP0_ipd, LGDEP0, VitalExtendToFillDelay(tipd_LGDEP0));
   VitalWireDelay (LGDEP1_ipd, LGDEP1, VitalExtendToFillDelay(tipd_LGDEP1));
   VitalWireDelay (LGDEP2_ipd, LGDEP2, VitalExtendToFillDelay(tipd_LGDEP2));
   VitalWireDelay (LEVEL0_ipd, LEVEL0, VitalExtendToFillDelay(tipd_LEVEL0));
   VitalWireDelay (LEVEL1_ipd, LEVEL1, VitalExtendToFillDelay(tipd_LEVEL1));
   VitalWireDelay (LEVEL2_ipd, LEVEL2, VitalExtendToFillDelay(tipd_LEVEL2));
   VitalWireDelay (LEVEL3_ipd, LEVEL3, VitalExtendToFillDelay(tipd_LEVEL3));
   VitalWireDelay (LEVEL4_ipd, LEVEL4, VitalExtendToFillDelay(tipd_LEVEL4));
   VitalWireDelay (LEVEL5_ipd, LEVEL5, VitalExtendToFillDelay(tipd_LEVEL5));
   VitalWireDelay (LEVEL6_ipd, LEVEL6, VitalExtendToFillDelay(tipd_LEVEL6));
   VitalWireDelay (LEVEL7_ipd, LEVEL7, VitalExtendToFillDelay(tipd_LEVEL7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RESET_ipd, RESET, VitalExtendToFillDelay(tipd_RESET));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (WCLKS_ipd, WCLKS, VitalExtendToFillDelay(tipd_WCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

   ---------------------------------------------------------------
   --                  Behavior Section                         --
   ---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);

    VITALBehavior : process (
                          LEVEL0_ipd, LEVEL1_ipd, LEVEL2_ipd, LEVEL3_ipd, LEVEL4_ipd, LEVEL5_ipd, LEVEL6_ipd, LEVEL7_ipd, 
                          LGDEP0_ipd, LGDEP1_ipd, LGDEP2_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd, RESET_ipd
                          )

     -- some internal veriable declaration
     variable RAM_di_int   : std_logic_vector(8 downto 0);
     variable memory_array : MEM_TYPE  := (others =>(others => 'X'));
     variable do_par       : std_logic := 'X';
     variable tmp_par      : std_logic := 'X';
     variable tmp_par2     : std_logic := 'X';
     variable wpe_var      : std_logic := 'X';
     variable temp         : integer   := 0;
     variable thresh       : integer   := 0;
     variable depth        : integer   := 0;
     variable WADDR        : integer   := 0;
     variable WADDR_wrap   : integer   := 0;
     variable RADDR        : integer   := 0;
     variable RADDR_wrap   : integer   := 0;

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     --  Read Timing Check Results
     variable PeriodData_RESET           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET                : X01                 := '0';
     variable Tviol_PARODD_RCLKS_posedge : X01                 := '0';
     variable TmDt_PARODD_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_RCLKS_posedge  : X01                 := '0';
     variable Tmkr_RESET_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable Tviol_DI0_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI0_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI1_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI2_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI3_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI4_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI5_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI6_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI7_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI8_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_PARODD_WCLKS_posedge : X01                 := '0';
     variable TmDt_PARODD_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_WCLKS_posedge    : X01                 := '0';
     variable TmDt_WRB_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_WCLKS_posedge  : X01                 := '0';
     variable TmDt_WBLKB_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_WCLKS_posedge  : X01                 := '0';
     variable Tmkr_RESET_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WCLKS                : X01                 := '0';

     -- functional Results


     variable DO0_zd   : std_ulogic;
     variable DO1_zd   : std_ulogic;
     variable DO2_zd   : std_ulogic;
     variable DO3_zd   : std_ulogic;
     variable DO4_zd   : std_ulogic;
     variable DO5_zd   : std_ulogic;
     variable DO6_zd   : std_ulogic;
     variable DO7_zd   : std_ulogic;
     variable DO8_zd   : std_ulogic;
     variable RPE_zd   : std_ulogic;
     variable WPE_zd   : std_ulogic;
     variable DOS_zd   : std_ulogic;
     variable FULL_zd  : std_ulogic;
     variable EMPTY_zd : std_ulogic;
     variable EQTH_zd  : std_ulogic;
     variable GEQTH_zd : std_ulogic;
     variable FULL_tmp  : std_ulogic;
     variable EMPTY_tmp : std_ulogic;
     variable EQTH_tmp  : std_ulogic;
     variable GEQTH_tmp : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData   : VitalGlitchDataType;
     variable DO1_GlitchData   : VitalGlitchDataType;
     variable DO2_GlitchData   : VitalGlitchDataType;
     variable DO3_GlitchData   : VitalGlitchDataType;
     variable DO4_GlitchData   : VitalGlitchDataType;
     variable DO5_GlitchData   : VitalGlitchDataType;
     variable DO6_GlitchData   : VitalGlitchDataType;
     variable DO7_GlitchData   : VitalGlitchDataType;
     variable DO8_GlitchData   : VitalGlitchDataType;
     variable RPE_GlitchData   : VitalGlitchDataType;
     variable WPE_GlitchData   : VitalGlitchDataType;
     variable DOS_GlitchData   : VitalGlitchDataType;
     variable FULL_GlitchData  : VitalGlitchDataType;
     variable EMPTY_GlitchData : VitalGlitchDataType;
     variable EQTH_GlitchData  : VitalGlitchDataType;
     variable GEQTH_GlitchData : VitalGlitchDataType;

     -- last value variables
     variable WCLKS_previous   : std_ulogic := 'X';
     variable RCLKS_previous   : std_ulogic := 'X';
     variable RBint_delayed    : std_ulogic := 'X';
     variable RBint_previous   : std_ulogic := 'X';
     variable WBint_delayed    : std_ulogic := 'X';
     variable WBint_previous   : std_ulogic := 'X';
     variable DIS_previous     : std_ulogic := 'X';
     variable RESET_previous   : std_ulogic := 'X';
     variable RESET_delayed    : std_ulogic := 'X';
     variable PARODD_previous  : std_ulogic := 'X';
     variable PARODD_delayed   : std_ulogic := 'X';
     variable DI0_delayed      : std_ulogic := 'X';
     variable DI1_delayed      : std_ulogic := 'X';
     variable DI2_delayed      : std_ulogic := 'X';
     variable DI3_delayed      : std_ulogic := 'X';
     variable DI4_delayed      : std_ulogic := 'X';
     variable DI5_delayed      : std_ulogic := 'X';
     variable DI6_delayed      : std_ulogic := 'X';
     variable DI7_delayed      : std_ulogic := 'X';
     variable DI8_delayed      : std_ulogic := 'X';
     variable DI0_previous     : std_ulogic := 'X';
     variable DI1_previous     : std_ulogic := 'X';
     variable DI2_previous     : std_ulogic := 'X';
     variable DI3_previous     : std_ulogic := 'X';
     variable DI4_previous     : std_ulogic := 'X';
     variable DI5_previous     : std_ulogic := 'X';
     variable DI6_previous     : std_ulogic := 'X';
     variable DI7_previous     : std_ulogic := 'X';
     variable DI8_previous     : std_ulogic := 'X';
     variable LGDEP0_delayed   : std_ulogic := 'X';
     variable LGDEP1_delayed   : std_ulogic := 'X';
     variable LGDEP2_delayed   : std_ulogic := 'X';
     variable LGDEP0_previous  : std_ulogic := 'X';
     variable LGDEP1_previous  : std_ulogic := 'X';
     variable LGDEP2_previous  : std_ulogic := 'X';
     variable LEVEL0_delayed   : std_ulogic := 'X';
     variable LEVEL1_delayed   : std_ulogic := 'X';
     variable LEVEL2_delayed   : std_ulogic := 'X';
     variable LEVEL3_delayed   : std_ulogic := 'X';
     variable LEVEL4_delayed   : std_ulogic := 'X';
     variable LEVEL5_delayed   : std_ulogic := 'X';
     variable LEVEL6_delayed   : std_ulogic := 'X';
     variable LEVEL7_delayed   : std_ulogic := 'X';
     variable LEVEL0_previous  : std_ulogic := 'X';
     variable LEVEL1_previous  : std_ulogic := 'X';
     variable LEVEL2_previous  : std_ulogic := 'X';
     variable LEVEL3_previous  : std_ulogic := 'X';
     variable LEVEL4_previous  : std_ulogic := 'X';
     variable LEVEL5_previous  : std_ulogic := 'X';
     variable LEVEL6_previous  : std_ulogic := 'X';
     variable LEVEL7_previous  : std_ulogic := 'X';

     -- Special variables to control flags
     variable hold_empty_low   : integer := 0;
     variable hold_eqth_high   : integer := 0;
     variable hold_geqth_high  : integer := 0;
     variable hold_full_low    : integer := 0;
     variable hold_empty_high  : integer := 0;
     variable hold_eqth_low    : integer := 0;
     variable hold_geqth_low   : integer := 0;

     variable WCLKS_re         : Time;
     variable WCLKS_fe         : Time;
     variable WCLKS_fe_prev    : Time;
     variable WB_re            : Time;
     variable RESET_re         : Time;


 begin -- process VITALBehavior

 if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

   -- recovery / removal check for RCLKS to RESET signal ;
       VitalRecoveryRemovalCheck ( Tviol_RESET_RCLKS_posedge,
                             Tmkr_RESET_RCLKS_posedge,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             trecovery_RESET_RCLKS_posedge_negedge,
                             thold_RESET_RCLKS_posedge_posedge,
                             TRUE,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'), 
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             TRUE,
                             TRUE,
                             WARNING
                             );

   -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             ((TO_X01(RBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             ((TO_X01(RDB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_PARODD_RCLKS_posedge,
                             TmDt_PARODD_RCLKS_posedge,
                             PARODD_ipd, "PARODD",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_PARODD_RCLKS_posedge_posedge,
                             tsetup_PARODD_RCLKS_negedge_posedge,
                             thold_PARODD_RCLKS_posedge_posedge,
                             thold_PARODD_RCLKS_negedge_posedge,
                             (TO_X01(RESET_ipd) = '1'),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (TO_X01(RDB) = '0') AND (TO_X01(RBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9SST",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RESET,
                              PeriodData_RESET,
                              RESET_ipd, "RESET",
                              0.0 ns,
                              tpw_RESET_negedge,
                              0.0 ns,
                              tpw_RESET_negedge,
                              True,
                              InstancePath & "/FIFO256x9SST",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       -- recovery / removal check for WCLKS to RESET signal ;
       VitalRecoveryRemovalCheck ( Tviol_RESET_WCLKS_posedge,
                             Tmkr_RESET_WCLKS_posedge,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns,
                             trecovery_RESET_WCLKS_posedge_negedge,
                             thold_RESET_WCLKS_posedge_posedge,
                             TRUE,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'), 
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             TRUE,
                             TRUE,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_posedge_posedge,
                             tsetup_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_posedge_posedge,
                             tsetup_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_posedge_posedge,
                             tsetup_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_posedge_posedge,
                             tsetup_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_posedge_posedge,
                             tsetup_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_posedge_posedge,
                             tsetup_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_posedge_posedge,
                             tsetup_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_posedge_posedge,
                             tsetup_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_posedge_posedge,
                             tsetup_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

   -- setup hold WEN, WBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_posedge_posedge,
                             tsetup_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_PARODD_WCLKS_posedge,
                             TmDt_PARODD_WCLKS_posedge,
                             PARODD_ipd, "PARODD",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_PARODD_WCLKS_posedge_posedge,
                             tsetup_PARODD_WCLKS_negedge_posedge,
                             thold_PARODD_WCLKS_posedge_posedge,
                             thold_PARODD_WCLKS_negedge_posedge,
                             ((TO_X01(RBint) = '0') AND (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/FIFO256x9SST",
                             True,
                             True,
                             WARNING
                             );

  --   Period of WCLK
      VitalPeriodPulseCheck ( Pviol_WCLKS,
                              PeriodData_WCLKS,
                              WCLKS_ipd, "WCLKS",
                              0.0 ns,
                              tperiod_WCLKS,
                              tpw_WCLKS_posedge,
                              tpw_WCLKS_negedge,
                              (TO_X01(WRB) = '0') AND (TO_X01(WBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9SST",
                              True,
                              True,
                              WARNING
                              );
 end if;

   ------------------------------------------------------------
   --               FIFO RESET                               --
   ------------------------------------------------------------

   if ( RESET_ipd'event and RESET_ipd = '0' ) then
       WADDR      := 0;
       RADDR      := 0;
       WADDR_wrap := 0;
       RADDR_wrap := 0;
       FULL_tmp   := '0';
       EMPTY_tmp  := '1';
       EQTH_tmp   := '0';
       GEQTH_tmp  := '0';
       WRITE_AT_PREV_EDGE <='0';
       READ_AT_PREV_EDGE <='0';
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
       hold_full_low   := 0;
       hold_empty_high := 0;
       hold_eqth_low   := 0;
       hold_geqth_low  := 0;
   end if;

   if ( WCLKS_ipd'event and WCLKS_ipd = '1' ) then
     WCLKS_re := now;
   end if;
      
   if ( WBint'event and WBint = '1' ) then
     WB_re := now;
   end if;
      
   if ( RESET_ipd'event and RESET_ipd = '1' ) then
     RESET_re := now;
     if ( TO_X01 ( WCLKS_ipd ) = '1' ) then
       if ( WCLKS_re = WB_re ) then
         hold_full_low   := 1; -- until next reset
         hold_empty_high := 1;
         hold_eqth_low   := 1;
         hold_geqth_low  := 1;
       elsif ( TO_X01 ( WBint ) = '0' ) then
         EMPTY_zd        := '0';
         EQTH_zd         := '1';
         GEQTH_zd        := '1';
         hold_empty_low  := 1; -- until next WCLKS falling edge
         hold_eqth_high  := 1;
         hold_geqth_high := 1;
       elsif ( WCLKS_re < WB_re ) then
         EMPTY_zd        := '0';
         EQTH_zd         := '1';
         GEQTH_zd        := '1';
         hold_empty_low  := 1; -- until next WCLKS falling edge
         hold_eqth_high  := 1;
         hold_geqth_high := 1;
       elsif ( WB_re < WCLKS_re ) then
         hold_empty_low  := 0; -- expected behavior
         hold_eqth_high  := 0;
         hold_geqth_high := 0;
         hold_full_low   := 0;
         hold_empty_high := 0;
         hold_eqth_low   := 0;
         hold_geqth_low  := 0;
       end if;
     else
       hold_empty_low  := 0; -- expected behavior
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
       hold_full_low   := 0;
       hold_empty_high := 0;
       hold_eqth_low   := 0;
       hold_geqth_low  := 0;
     end if;
   end if;

   if ( WCLKS_ipd'event and WCLKS_ipd = '0' ) then
     WCLKS_fe_prev := WCLKS_fe;
     WCLKS_fe := now;
     if (( TO_X01 ( RESET_ipd ) = '1' ) and ( WCLKS_fe_prev < RESET_re )) then
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
     end if;
   end if;


   ------------------------------------------------------------
   --    wpe output                                           -
   ------------------------------------------------------------

   if ( PARODD_ipd'EVENT ) then
     RPE_zd   := not RPE_zd;
     WPE_zd := not WPE_zd;
   end if;

   ------------------------------------------------------------
   --         WPE generating block                            -
   ------------------------------------------------------------

    if (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
        tmp_par := DI7_delayed XOR DI6_delayed XOR DI5_delayed XOR DI4_delayed XOR DI3_delayed XOR DI2_delayed XOR DI1_delayed XOR DI0_delayed;
        par_f    <= tmp_par ;
        tmp_par2 := (tmp_par xor DI8_delayed);
        par_f2   <= tmp_par2;

      if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
          ( TO_X01 ( DI8_ipd )    = 'X' ) or
          ( TO_X01 ( DI7_ipd )    = 'X' ) or
          ( TO_X01 ( DI6_ipd )    = 'X' ) or
          ( TO_X01 ( DI5_ipd )    = 'X' ) or
          ( TO_X01 ( DI4_ipd )    = 'X' ) or
          ( TO_X01 ( DI3_ipd )    = 'X' ) or
          ( TO_X01 ( DI2_ipd )    = 'X' ) or
          ( TO_X01 ( DI1_ipd )    = 'X' ) or
          ( TO_X01 ( DI0_ipd )    = 'X' )
         ) then
        wpe_var  :=  'X';
      else
        if ( tmp_par2 /= PARODD_ipd ) then
          wpe_var  :=  '1';
        else
          wpe_var  :=  '0';
        end if;
      end if;
        RAM_di_int(8) := DI8_delayed;
        WPE_zd := wpe_var;
    end if;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

   if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
   end if; 

   -----------------------------------------------------------
   --    calculate the depth and levels                     --
   -----------------------------------------------------------

    temp :=((INT(LGDEP2_delayed)*4) + (INT(LGDEP1_delayed)*2) + 
           (INT(LGDEP0_delayed)*1));

    case temp is 
         when 0 => depth := 2;
         when 1 => depth := 4;
         when 2 => depth := 8;
         when 3 => depth := 16;
         when 4 => depth := 32;
         when 5 => depth := 64;
         when 6 => depth := 128;
         when 7 => depth := 256;
         when others => depth := 0;
    end case;

    -- thresh value

    thresh := (INT(LEVEL7_delayed)*128) + (INT(LEVEL6_delayed)*64) + 
               (INT(LEVEL5_delayed)*32) + (INT(LEVEL4_delayed)*16) + 
               (INT(LEVEL3_delayed)*8) + (INT(LEVEL2_delayed)*4) + 
               (INT(LEVEL1_delayed)*2) + (INT(LEVEL0_delayed)*1); 

    if ( thresh = 0 or thresh = 255 ) then
      assert false
        report " Illegal level configuration, LEVEL cannot be 0 or 255 "
        severity failure;
    end if;

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

   if(TO_X01(WCLKS_ipd)='X') then
    if(RESET_delayed = '1') then
     if (WBint_delayed = '0') then
      if (TO_X01(WCLKS_previous) /= 'X') then
        assert false
        report ": WCLK unknown"
        severity Error;
      end if;
     end if;
    end if;
   elsif (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') AND (TO_X01(RESET_ipd) = '1')then
     WRITE_AT_PREV_EDGE <='0';
     case (TO_X01(WBint_delayed)) is 
      when '1' =>
                null;
      when '0' => 
         if(FULL_zd = '0') then 
         RAM_di_int(7 downto 0) := DI7_delayed & DI6_delayed & DI5_delayed & 
                                    DI4_delayed & DI3_delayed & DI2_delayed & 
                                    DI1_delayed & DI0_delayed;
         memory_array(WADDR) := RAM_di_int;
         WRITE_AT_PREV_EDGE <='1';
         if(WADDR <depth-1  ) then
           WADDR := WADDR + 1;
         elsif( WADDR  = depth-1) then
           WADDR := 0;
           WADDR_wrap := 1 - WADDR_wrap;
         end if;
        end if;
       when others => 
        if (TO_X01(WBint_previous) /= 'X') then
          assert false
          report ": WBLKB or WRB unknown"
          severity Error;
          end if;
        end case;
     elsif(WCLKS_ipd'EVENT AND WCLKS_ipd = '0')  AND (TO_X01(RESET_delayed) = '1') AND (TO_X01(WRITE_AT_PREV_EDGE) = '1')then
        WRITE_AT_PREV_EDGE <='0';
        if(WADDR   = RADDR ) then
         if(RADDR_wrap /= WADDR_wrap) then
          FULL_tmp := '1';
          EMPTY_tmp :='0';
         end if;
        end if;
        if(WADDR   /= RADDR ) then
          EMPTY_tmp := '0';
        end if;
          if(RADDR_wrap = WADDR_wrap) then
            if(WADDR - RADDR = thresh ) then
               EQTH_tmp := '1';
            else 
               EQTH_tmp := '0';
            end if;
            if(WADDR - RADDR >= thresh ) then
                GEQTH_tmp := '1';
            else 
                GEQTH_tmp := '0';
            end if;
          else 
           if((depth -RADDR + WADDR) = thresh ) then
               EQTH_tmp := '1';
            else 
               EQTH_tmp := '0';
            end if;
            if((depth -RADDR + WADDR) >= thresh ) then
                GEQTH_tmp := '1';
            else 
                GEQTH_tmp := '0';
            end if;
           end if; 
      else
       null;
    end if;


  --------------------------------------------------------------------
  --          FIFO READ SECTION........                             --
  --------------------------------------------------------------------

  if (TO_X01(RCLKS_ipd)='X') then
    if(RESET_ipd /= '0') then
    if(TO_X01(RBint_delayed) /= '1') then
      if(TO_X01(RCLKS_previous) /= 'X') then
        assert false
        report ": RCLK unknown"
        severity Error;
        DO0_zd  := 'X';
        DO1_zd  := 'X';
        DO2_zd  := 'X';
        DO3_zd  := 'X';
        DO4_zd  := 'X';
        DO5_zd  := 'X';
        DO6_zd  := 'X';
        DO7_zd  := 'X';
        DO8_zd  := 'X';
      end if;
     end if;
    end if;
   elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='1') AND (TO_X01(RESET_delayed) = '1')) then
     READ_AT_PREV_EDGE <='0';
     case (TO_X01(RBint_delayed)) is
        when '1' =>
                null;
        when '0' =>
         if(TO_X01(EMPTY_zd) /= '1') then 
           DO0_zd  := memory_array(RADDR)(0);
           DO1_zd  := memory_array(RADDR)(1);
           DO2_zd  := memory_array(RADDR)(2);
           DO3_zd  := memory_array(RADDR)(3);
           DO4_zd  := memory_array(RADDR)(4);
           DO5_zd  := memory_array(RADDR)(5);
           DO6_zd  := memory_array(RADDR)(6);
           DO7_zd  := memory_array(RADDR)(7);
           DO8_zd  := memory_array(RADDR)(8);
           READ_AT_PREV_EDGE <='1';
           if(RADDR <depth-1  ) then
             RADDR := RADDR + 1;
           else
             RADDR :=(RADDR +1) mod  depth;
             RADDR_wrap :=1 - RADDR_wrap;
           end if;
            do_par  := DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR DO3_zd XOR
                       DO2_zd XOR DO1_zd XOR DO0_zd;
            par_f <= do_par;
            if (do_par = 'X') then
             RPE_zd := 'X';
            elsif (do_par /= PARODD_delayed) then
             RPE_zd  :=  '1';
            else
             RPE_zd  :=  '0';
            end if;
         end if;
     when others =>
       if (TO_X01(RBint_previous) /= 'X') then
        assert false
        report ": RDB or RBLKB unknown"
        severity Error;
        end if;
           DO0_zd  := 'X';
           DO1_zd  := 'X';
           DO2_zd  := 'X';
           DO3_zd  := 'X';
           DO4_zd  := 'X';
           DO5_zd  := 'X';
           DO6_zd  := 'X';
           DO7_zd  := 'X';
           DO8_zd  := 'X';
     end case;
  elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='0') AND (TO_X01(RESET_delayed) = '1') AND (TO_X01(READ_AT_PREV_EDGE) = '1')) then
   READ_AT_PREV_EDGE <='0';
   if(RADDR = WADDR ) then
    if(RADDR_wrap = WADDR_wrap) then
       EMPTY_tmp := '1';
       FULL_tmp  := '0';
    end if;
   end if;
   if(RADDR /= WADDR ) then
    FULL_tmp  := '0';
   end if;
    if(WADDR_wrap = RADDR_wrap ) then
     if((WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((WADDR - RADDR) >= thresh  ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    else 
     if((depth + WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((depth + WADDR - RADDR) >= thresh ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    end if;
 else 
    null;
 end if;

   -- Mimic odd silicon flag behavior coming out of RESET with WB low
   
   if ( hold_full_low = 1 ) then
     FULL_zd := '0';
   else
     FULL_zd := FULL_tmp;
   end if;

   if ( hold_empty_low = 1 ) then
     EMPTY_zd := '0';
   elsif ( hold_empty_high = 1 ) then
     EMPTY_zd := '1';
   else
     EMPTY_zd := EMPTY_tmp;
   end if;

   if ( hold_eqth_high = 1 ) then
     EQTH_zd := '1';
   elsif ( hold_eqth_low = 1 ) then
     EQTH_zd := '0';
   else
     EQTH_zd := EQTH_tmp;
   end if;

   -- If LEVEL greater than DEPTH then GEQTH mimics FULL
   
   if ( hold_geqth_high = 1 ) then
     GEQTH_zd := '1';
   elsif ( hold_geqth_low = 1 ) then
     GEQTH_zd := '0';
   else
     if ( thresh > depth ) then
       GEQTH_zd := FULL_zd;
     else
       GEQTH_zd := GEQTH_tmp;
     end if;
   end if;


  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       WCLKS_previous  := WCLKS_ipd;
       RCLKS_previous   := RCLKS_ipd;
       RBint_previous   := RBint_delayed;
       RBint_delayed    := RBint;
       WBint_previous   := WBint_delayed;
       WBint_delayed    := WBint;
       DI0_delayed      := DI0_ipd;
       DI1_delayed      := DI1_ipd;
       DI2_delayed      := DI2_ipd;
       DI3_delayed      := DI3_ipd;
       DI4_delayed      := DI4_ipd;
       DI5_delayed      := DI5_ipd;
       DI6_delayed      := DI6_ipd;
       DI7_delayed      := DI7_ipd;
       DI8_delayed      := DI8_ipd;
       LGDEP0_previous  := LGDEP0_delayed;
       LGDEP0_delayed   := LGDEP0_ipd;
       LGDEP1_previous  := LGDEP1_delayed;
       LGDEP1_delayed   := LGDEP1_ipd;
       LGDEP2_previous  := LGDEP2_delayed;
       LGDEP2_delayed   := LGDEP2_ipd;
       LEVEL0_previous  := LEVEL0_delayed;
       LEVEL0_delayed   := LEVEL0_ipd;
       LEVEL1_previous  := LEVEL1_delayed;
       LEVEL1_delayed   := LEVEL1_ipd;
       LEVEL2_previous  := LEVEL2_delayed;
       LEVEL2_delayed   := LEVEL2_ipd;
       LEVEL3_previous  := LEVEL3_delayed;
       LEVEL3_delayed   := LEVEL3_ipd;
       LEVEL4_previous  := LEVEL4_delayed;
       LEVEL4_delayed   := LEVEL4_ipd;
       LEVEL5_previous  := LEVEL5_delayed;
       LEVEL5_delayed   := LEVEL5_ipd;
       LEVEL6_previous  := LEVEL6_delayed;
       LEVEL6_delayed   := LEVEL6_ipd;
       LEVEL7_previous  := LEVEL7_delayed;
       LEVEL7_delayed   := LEVEL7_ipd;
       PARODD_previous  := PARODD_delayed; 
       PARODD_delayed   := PARODD_ipd;
       RESET_previous   := RESET_delayed; 
       RESET_delayed    := RESET_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
             OutSignal     => DOS,
             GlitchData    => DOS_GlitchData,
             OutSignalName => "DOS",
             OutTemp       => DOS_zd,

             Paths =>   (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
           OutSignal     => WPE,
           GlitchData    => WPE_GlitchData,
           OutSignalName => "WPE",
           OutTemp       => WPE_zd,
           Paths =>   (0  => (WCLKS_ipd'last_event,
                       VitalExtendToFillDelay(tpd_WCLKS_WPE), true),
                       1 => (PARODD_ipd'last_event,
                             VitalExtendToFillDelay(tpd_PARODD_WPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO0), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO1), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO2), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO3), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO4), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO5), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO6), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO7), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO8), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => RPE,
           GlitchData    => RPE_GlitchData,
           OutSignalName => "RPE",
           OutTemp       => RPE_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_RPE), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_RPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => FULL,
           GlitchData    => FULL_GlitchData,
           OutSignalName => "FULL",
           OutTemp       => FULL_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_FULL), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_FULL), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_FULL), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EMPTY,
           GlitchData    => EMPTY_GlitchData,
           OutSignalName => "EMPTY",
           OutTemp       => EMPTY_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EMPTY), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_EMPTY), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EMPTY), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EQTH,
           GlitchData    => EQTH_GlitchData,
           OutSignalName => "EQTH",
           OutTemp       => EQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EQTH), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_EQTH), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => GEQTH,
           GlitchData    => GEQTH_GlitchData,
           OutSignalName => "GEQTH",
           OutTemp       => GEQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_GEQTH), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_GEQTH), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_GEQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );


   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

LIBRARY a500k;
USE a500k.all;

entity FIFO256x9SSTP is 
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_WCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_WCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;

        -- WCLK falling edge setup to RESET rising edge 
 	trecovery_RESET_WCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_WCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- WCLK rising  edge hold to RESET rising edge 
	thold_RESET_WCLKS_posedge_posedge             : VitalDelayType := 0.00 ns;
	thold_RESET_WCLKS_posedge_negedge             : VitalDelayType := 0.00 ns;
	tpw_WCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        WCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');


ATTRIBUTE VITAL_LEVEL0 OF FIFO256x9SSTP : entity IS True ;
END FIFO256x9SSTP;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of FIFO256x9SSTP is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal LGDEP0_ipd : std_ulogic := 'X';
   signal LGDEP1_ipd : std_ulogic := 'X';
   signal LGDEP2_ipd : std_ulogic := 'X';
   signal LEVEL0_ipd : std_ulogic := 'X';
   signal LEVEL1_ipd : std_ulogic := 'X';
   signal LEVEL2_ipd : std_ulogic := 'X';
   signal LEVEL3_ipd : std_ulogic := 'X';
   signal LEVEL4_ipd : std_ulogic := 'X';
   signal LEVEL5_ipd : std_ulogic := 'X';
   signal LEVEL6_ipd : std_ulogic := 'X';
   signal LEVEL7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal RESET_ipd  : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal WCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

   -- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic := 'X';
   signal par_f2     : std_logic := 'X';

   signal WRITE_AT_PREV_EDGE : std_logic := '0';
   signal READ_AT_PREV_EDGE  : std_logic := '0';

   begin  --  VITAL_ACT

   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (LGDEP0_ipd, LGDEP0, VitalExtendToFillDelay(tipd_LGDEP0));
   VitalWireDelay (LGDEP1_ipd, LGDEP1, VitalExtendToFillDelay(tipd_LGDEP1));
   VitalWireDelay (LGDEP2_ipd, LGDEP2, VitalExtendToFillDelay(tipd_LGDEP2));
   VitalWireDelay (LEVEL0_ipd, LEVEL0, VitalExtendToFillDelay(tipd_LEVEL0));
   VitalWireDelay (LEVEL1_ipd, LEVEL1, VitalExtendToFillDelay(tipd_LEVEL1));
   VitalWireDelay (LEVEL2_ipd, LEVEL2, VitalExtendToFillDelay(tipd_LEVEL2));
   VitalWireDelay (LEVEL3_ipd, LEVEL3, VitalExtendToFillDelay(tipd_LEVEL3));
   VitalWireDelay (LEVEL4_ipd, LEVEL4, VitalExtendToFillDelay(tipd_LEVEL4));
   VitalWireDelay (LEVEL5_ipd, LEVEL5, VitalExtendToFillDelay(tipd_LEVEL5));
   VitalWireDelay (LEVEL6_ipd, LEVEL6, VitalExtendToFillDelay(tipd_LEVEL6));
   VitalWireDelay (LEVEL7_ipd, LEVEL7, VitalExtendToFillDelay(tipd_LEVEL7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RESET_ipd, RESET, VitalExtendToFillDelay(tipd_RESET));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (WCLKS_ipd, WCLKS, VitalExtendToFillDelay(tipd_WCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

   ---------------------------------------------------------------
   --                  Behavior Section                         --
   ---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);

    VITALBehavior : process (
                          LEVEL0_ipd, LEVEL1_ipd, LEVEL2_ipd, LEVEL3_ipd, LEVEL4_ipd, LEVEL5_ipd, LEVEL6_ipd, LEVEL7_ipd, 
                          LGDEP0_ipd, LGDEP1_ipd, LGDEP2_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd, RESET_ipd
                          )

     -- some internal veriable declaration
     variable RAM_di_int   : std_logic_vector(8 downto 0);
     variable memory_array : MEM_TYPE  := (others =>(others => 'X'));
     variable do_par       : std_logic := 'X';
     variable tmp_par      : std_logic := 'X';
     variable tmp_par2     : std_logic := 'X';
     variable wpe_var      : std_logic := 'X';
     variable temp         : integer   := 0;
     variable thresh       : integer   := 0;
     variable depth        : integer   := 0;
     variable WADDR        : integer   := 0;
     variable WADDR_wrap   : integer   := 0;
     variable RADDR        : integer   := 0;
     variable RADDR_wrap   : integer   := 0;

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     --  Read Timing Check Results
     variable PeriodData_RESET           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET                : X01                 := '0';
     variable Tviol_PARODD_RCLKS_posedge : X01                 := '0';
     variable TmDt_PARODD_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_RCLKS_posedge  : X01                 := '0';
     variable Tmkr_RESET_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable Tviol_DI0_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI0_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI1_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI2_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI3_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI4_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI5_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI6_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI7_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI8_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_PARODD_WCLKS_posedge : X01                 := '0';
     variable TmDt_PARODD_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_WCLKS_posedge    : X01                 := '0';
     variable TmDt_WRB_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_WCLKS_posedge  : X01                 := '0';
     variable TmDt_WBLKB_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_WCLKS_posedge  : X01                 := '0';
     variable Tmkr_RESET_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WCLKS                : X01                 := '0';

     -- functional Results


     variable DO0_zd   : std_ulogic;
     variable DO1_zd   : std_ulogic;
     variable DO2_zd   : std_ulogic;
     variable DO3_zd   : std_ulogic;
     variable DO4_zd   : std_ulogic;
     variable DO5_zd   : std_ulogic;
     variable DO6_zd   : std_ulogic;
     variable DO7_zd   : std_ulogic;
     variable DO8_zd   : std_ulogic;
     variable RPE_zd   : std_ulogic;
     variable WPE_zd   : std_ulogic;
     variable DOS_zd   : std_ulogic;
     variable FULL_zd  : std_ulogic;
     variable EMPTY_zd : std_ulogic;
     variable EQTH_zd  : std_ulogic;
     variable GEQTH_zd : std_ulogic;
     variable FULL_tmp  : std_ulogic;
     variable EMPTY_tmp : std_ulogic;
     variable EQTH_tmp  : std_ulogic;
     variable GEQTH_tmp : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData   : VitalGlitchDataType;
     variable DO1_GlitchData   : VitalGlitchDataType;
     variable DO2_GlitchData   : VitalGlitchDataType;
     variable DO3_GlitchData   : VitalGlitchDataType;
     variable DO4_GlitchData   : VitalGlitchDataType;
     variable DO5_GlitchData   : VitalGlitchDataType;
     variable DO6_GlitchData   : VitalGlitchDataType;
     variable DO7_GlitchData   : VitalGlitchDataType;
     variable DO8_GlitchData   : VitalGlitchDataType;
     variable DOS_GlitchData   : VitalGlitchDataType;
     variable FULL_GlitchData  : VitalGlitchDataType;
     variable EMPTY_GlitchData : VitalGlitchDataType;
     variable EQTH_GlitchData  : VitalGlitchDataType;
     variable GEQTH_GlitchData : VitalGlitchDataType;

     -- last value variables
     variable WCLKS_previous   : std_ulogic := 'X';
     variable RCLKS_previous   : std_ulogic := 'X';
     variable RBint_delayed    : std_ulogic := 'X';
     variable RBint_previous   : std_ulogic := 'X';
     variable WBint_delayed    : std_ulogic := 'X';
     variable WBint_previous   : std_ulogic := 'X';
     variable DIS_previous     : std_ulogic := 'X';
     variable RESET_previous   : std_ulogic := 'X';
     variable RESET_delayed    : std_ulogic := 'X';
     variable PARODD_previous  : std_ulogic := 'X';
     variable PARODD_delayed   : std_ulogic := 'X';
     variable DI0_delayed      : std_ulogic := 'X';
     variable DI1_delayed      : std_ulogic := 'X';
     variable DI2_delayed      : std_ulogic := 'X';
     variable DI3_delayed      : std_ulogic := 'X';
     variable DI4_delayed      : std_ulogic := 'X';
     variable DI5_delayed      : std_ulogic := 'X';
     variable DI6_delayed      : std_ulogic := 'X';
     variable DI7_delayed      : std_ulogic := 'X';
     variable DI8_delayed      : std_ulogic := 'X';
     variable DI0_previous     : std_ulogic := 'X';
     variable DI1_previous     : std_ulogic := 'X';
     variable DI2_previous     : std_ulogic := 'X';
     variable DI3_previous     : std_ulogic := 'X';
     variable DI4_previous     : std_ulogic := 'X';
     variable DI5_previous     : std_ulogic := 'X';
     variable DI6_previous     : std_ulogic := 'X';
     variable DI7_previous     : std_ulogic := 'X';
     variable DI8_previous     : std_ulogic := 'X';
     variable LGDEP0_delayed   : std_ulogic := 'X';
     variable LGDEP1_delayed   : std_ulogic := 'X';
     variable LGDEP2_delayed   : std_ulogic := 'X';
     variable LGDEP0_previous  : std_ulogic := 'X';
     variable LGDEP1_previous  : std_ulogic := 'X';
     variable LGDEP2_previous  : std_ulogic := 'X';
     variable LEVEL0_delayed   : std_ulogic := 'X';
     variable LEVEL1_delayed   : std_ulogic := 'X';
     variable LEVEL2_delayed   : std_ulogic := 'X';
     variable LEVEL3_delayed   : std_ulogic := 'X';
     variable LEVEL4_delayed   : std_ulogic := 'X';
     variable LEVEL5_delayed   : std_ulogic := 'X';
     variable LEVEL6_delayed   : std_ulogic := 'X';
     variable LEVEL7_delayed   : std_ulogic := 'X';
     variable LEVEL0_previous  : std_ulogic := 'X';
     variable LEVEL1_previous  : std_ulogic := 'X';
     variable LEVEL2_previous  : std_ulogic := 'X';
     variable LEVEL3_previous  : std_ulogic := 'X';
     variable LEVEL4_previous  : std_ulogic := 'X';
     variable LEVEL5_previous  : std_ulogic := 'X';
     variable LEVEL6_previous  : std_ulogic := 'X';
     variable LEVEL7_previous  : std_ulogic := 'X';

     -- Special variables to control flags
     variable hold_empty_low   : integer := 0;
     variable hold_eqth_high   : integer := 0;
     variable hold_geqth_high  : integer := 0;
     variable hold_full_low    : integer := 0;
     variable hold_empty_high  : integer := 0;
     variable hold_eqth_low    : integer := 0;
     variable hold_geqth_low   : integer := 0;

     variable WCLKS_re         : Time;
     variable WCLKS_fe         : Time;
     variable WCLKS_fe_prev    : Time;
     variable WB_re            : Time;
     variable RESET_re         : Time;


 begin -- process VITALBehavior

 if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

   -- recovery / removal check for RCLKS to RESET signal ;
       VitalRecoveryRemovalCheck ( Tviol_RESET_RCLKS_posedge,
                             Tmkr_RESET_RCLKS_posedge,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             trecovery_RESET_RCLKS_posedge_negedge,
                             thold_RESET_RCLKS_posedge_posedge,
                             TRUE,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'), 
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             TRUE,
                             TRUE,
                             WARNING
                             );

   -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             ((TO_X01(RBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             ((TO_X01(RDB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_PARODD_RCLKS_posedge,
                             TmDt_PARODD_RCLKS_posedge,
                             PARODD_ipd, "PARODD",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_PARODD_RCLKS_posedge_posedge,
                             tsetup_PARODD_RCLKS_negedge_posedge,
                             thold_PARODD_RCLKS_posedge_posedge,
                             thold_PARODD_RCLKS_negedge_posedge,
                             (TO_X01(RESET_ipd) = '1'),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (TO_X01(RDB) = '0') AND (TO_X01(RBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9SSTP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RESET,
                              PeriodData_RESET,
                              RESET_ipd, "RESET",
                              0.0 ns,
                              tpw_RESET_negedge,
                              0.0 ns,
                              tpw_RESET_negedge,
                              True,
                              InstancePath & "/FIFO256x9SSTP",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       -- recovery / removal check for WCLKS to RESET signal ;
       VitalRecoveryRemovalCheck ( Tviol_RESET_WCLKS_posedge,
                             Tmkr_RESET_WCLKS_posedge,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns,
                             trecovery_RESET_WCLKS_posedge_negedge,
                             thold_RESET_WCLKS_posedge_posedge,
                             TRUE,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'), 
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             TRUE,
                             TRUE,
                             WARNING
                             );

       -- setup /hold check for WCLK to RESET signal ;
       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_posedge_posedge,
                             tsetup_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_posedge_posedge,
                             tsetup_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_posedge_posedge,
                             tsetup_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_posedge_posedge,
                             tsetup_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_posedge_posedge,
                             tsetup_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_posedge_posedge,
                             tsetup_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_posedge_posedge,
                             tsetup_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_posedge_posedge,
                             tsetup_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_posedge_posedge,
                             tsetup_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

   -- setup hold WEN, WBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_posedge_posedge,
                             tsetup_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_PARODD_WCLKS_posedge,
                             TmDt_PARODD_WCLKS_posedge,
                             PARODD_ipd, "PARODD",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_PARODD_WCLKS_posedge_posedge,
                             tsetup_PARODD_WCLKS_negedge_posedge,
                             thold_PARODD_WCLKS_posedge_posedge,
                             thold_PARODD_WCLKS_negedge_posedge,
                             ((TO_X01(RBint) = '0') AND (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/FIFO256x9SSTP",
                             True,
                             True,
                             WARNING
                             );

  --   Period of WCLK
      VitalPeriodPulseCheck ( Pviol_WCLKS,
                              PeriodData_WCLKS,
                              WCLKS_ipd, "WCLKS",
                              0.0 ns,
                              tperiod_WCLKS,
                              tpw_WCLKS_posedge,
                              tpw_WCLKS_negedge,
                              (TO_X01(WRB) = '0') AND (TO_X01(WBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9SSTP",
                              True,
                              True,
                              WARNING
                              );
 end if;

   ------------------------------------------------------------
   --               FIFO RESET                               --
   ------------------------------------------------------------

   if ( RESET_ipd'event and RESET_ipd = '0' ) then
       WADDR      := 0;
       RADDR      := 0;
       WADDR_wrap := 0;
       RADDR_wrap := 0;
       FULL_tmp   := '0';
       EMPTY_tmp  := '1';
       EQTH_tmp   := '0';
       GEQTH_tmp  := '0';
       WRITE_AT_PREV_EDGE <='0';
       READ_AT_PREV_EDGE <='0';
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
       hold_full_low   := 0;
       hold_empty_high := 0;
       hold_eqth_low   := 0;
       hold_geqth_low  := 0;
   end if;

   if ( WCLKS_ipd'event and WCLKS_ipd = '1' ) then
     WCLKS_re := now;
   end if;
      
   if ( WBint'event and WBint = '1' ) then
     WB_re := now;
   end if;
      
   if ( RESET_ipd'event and RESET_ipd = '1' ) then
     RESET_re := now;
     if ( TO_X01 ( WCLKS_ipd ) = '1' ) then
       if ( WCLKS_re = WB_re ) then
         hold_full_low   := 1; -- until next reset
         hold_empty_high := 1;
         hold_eqth_low   := 1;
         hold_geqth_low  := 1;
       elsif ( TO_X01 ( WBint ) = '0' ) then
         EMPTY_zd        := '0';
         EQTH_zd         := '1';
         GEQTH_zd        := '1';
         hold_empty_low  := 1; -- until next WCLKS falling edge
         hold_eqth_high  := 1;
         hold_geqth_high := 1;
       elsif ( WCLKS_re < WB_re ) then
         EMPTY_zd        := '0';
         EQTH_zd         := '1';
         GEQTH_zd        := '1';
         hold_empty_low  := 1; -- until next WCLKS falling edge
         hold_eqth_high  := 1;
         hold_geqth_high := 1;
       elsif ( WB_re < WCLKS_re ) then
         hold_empty_low  := 0; -- expected behavior
         hold_eqth_high  := 0;
         hold_geqth_high := 0;
         hold_full_low   := 0;
         hold_empty_high := 0;
         hold_eqth_low   := 0;
         hold_geqth_low  := 0;
       end if;
     else
       hold_empty_low  := 0; -- expected behavior
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
       hold_full_low   := 0;
       hold_empty_high := 0;
       hold_eqth_low   := 0;
       hold_geqth_low  := 0;
     end if;
   end if;

   if ( WCLKS_ipd'event and WCLKS_ipd = '0' ) then
     WCLKS_fe_prev := WCLKS_fe;
     WCLKS_fe := now;
     if (( TO_X01 ( RESET_ipd ) = '1' ) and ( WCLKS_fe_prev < RESET_re )) then
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
     end if;
   end if;


   ------------------------------------------------------------
   --         WPE generating block                            -
   ------------------------------------------------------------

    if (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      tmp_par  := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;
      par_f  <= tmp_par ;
      if (tmp_par /= PARODD_ipd) then
        wpe_var  :=  '1';
      else
        wpe_var  :=  '0';
      end if;
      RAM_di_int(8) := wpe_var;
      WPE_zd := wpe_var;
    end if;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

   if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
   end if; 

   -----------------------------------------------------------
   --    calculate the depth and levels                     --
   -----------------------------------------------------------

    temp :=((INT(LGDEP2_delayed)*4) + (INT(LGDEP1_delayed)*2) + 
           (INT(LGDEP0_delayed)*1));

    case temp is 
         when 0 => depth := 2;
         when 1 => depth := 4;
         when 2 => depth := 8;
         when 3 => depth := 16;
         when 4 => depth := 32;
         when 5 => depth := 64;
         when 6 => depth := 128;
         when 7 => depth := 256;
         when others => depth := 0;
    end case;

    -- thresh value

    thresh := (INT(LEVEL7_delayed)*128) + (INT(LEVEL6_delayed)*64) + 
               (INT(LEVEL5_delayed)*32) + (INT(LEVEL4_delayed)*16) + 
               (INT(LEVEL3_delayed)*8) + (INT(LEVEL2_delayed)*4) + 
               (INT(LEVEL1_delayed)*2) + (INT(LEVEL0_delayed)*1); 

    if ( thresh = 0 or thresh = 255 ) then
      assert false
        report " Illegal level configuration, LEVEL cannot be 0 or 255 "
        severity failure;
    end if;

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

   if(TO_X01(WCLKS_ipd)='X') then
    if(RESET_delayed = '1') then
     if (WBint_delayed = '0') then
      if (TO_X01(WCLKS_previous) /= 'X') then
        assert false
        report ": WCLK unknown"
        severity Error;
      end if;
     end if;
    end if;
   elsif (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') AND (TO_X01(RESET_ipd) = '1')then
     WRITE_AT_PREV_EDGE <='0';
     case (TO_X01(WBint_delayed)) is 
      when '1' =>
                null;
      when '0' => 
         if(FULL_zd = '0') then 
         RAM_di_int(7 downto 0) := DI7_delayed & DI6_delayed & DI5_delayed & 
                                    DI4_delayed & DI3_delayed & DI2_delayed & 
                                    DI1_delayed & DI0_delayed;
         memory_array(WADDR) := RAM_di_int;
         WRITE_AT_PREV_EDGE <='1';
         if(WADDR <depth-1  ) then
           WADDR := WADDR + 1;
         elsif( WADDR  = depth-1) then
           WADDR := 0;
           WADDR_wrap := 1 - WADDR_wrap;
         end if;
        end if;
       when others => 
        if (TO_X01(WBint_previous) /= 'X') then
          assert false
          report ": WBLKB or WRB unknown"
          severity Error;
          end if;
        end case;
     elsif(WCLKS_ipd'EVENT AND WCLKS_ipd = '0')  AND (TO_X01(RESET_delayed) = '1') AND (TO_X01(WRITE_AT_PREV_EDGE) = '1')then
        WRITE_AT_PREV_EDGE <='0';
        if(WADDR   = RADDR ) then
         if(RADDR_wrap /= WADDR_wrap) then
          FULL_tmp := '1';
          EMPTY_tmp :='0';
         end if;
        end if;
        if(WADDR   /= RADDR ) then
          EMPTY_tmp := '0';
        end if;
          if(RADDR_wrap = WADDR_wrap) then
            if(WADDR - RADDR = thresh ) then
               EQTH_tmp := '1';
            else 
               EQTH_tmp := '0';
            end if;
            if(WADDR - RADDR >= thresh ) then
                GEQTH_tmp := '1';
            else 
                GEQTH_tmp := '0';
            end if;
          else 
           if((depth -RADDR + WADDR) = thresh ) then
               EQTH_tmp := '1';
            else 
               EQTH_tmp := '0';
            end if;
            if((depth -RADDR + WADDR) >= thresh ) then
                GEQTH_tmp := '1';
            else 
                GEQTH_tmp := '0';
            end if;
           end if; 
      else
       null;
    end if;


  --------------------------------------------------------------------
  --          FIFO READ SECTION........                             --
  --------------------------------------------------------------------

  if (TO_X01(RCLKS_ipd)='X') then
    if(RESET_ipd /= '0') then
    if(TO_X01(RBint_delayed) /= '1') then
      if(TO_X01(RCLKS_previous) /= 'X') then
        assert false
        report ": RCLK unknown"
        severity Error;
        DO0_zd  := 'X';
        DO1_zd  := 'X';
        DO2_zd  := 'X';
        DO3_zd  := 'X';
        DO4_zd  := 'X';
        DO5_zd  := 'X';
        DO6_zd  := 'X';
        DO7_zd  := 'X';
        DO8_zd  := 'X';
      end if;
     end if;
    end if;
   elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='1') AND (TO_X01(RESET_delayed) = '1')) then
     READ_AT_PREV_EDGE <='0';
     case (TO_X01(RBint_delayed)) is
        when '1' =>
                null;
        when '0' =>
         if(TO_X01(EMPTY_zd) /= '1') then 
           DO0_zd  := memory_array(RADDR)(0);
           DO1_zd  := memory_array(RADDR)(1);
           DO2_zd  := memory_array(RADDR)(2);
           DO3_zd  := memory_array(RADDR)(3);
           DO4_zd  := memory_array(RADDR)(4);
           DO5_zd  := memory_array(RADDR)(5);
           DO6_zd  := memory_array(RADDR)(6);
           DO7_zd  := memory_array(RADDR)(7);
           DO8_zd  := memory_array(RADDR)(8);
           READ_AT_PREV_EDGE <='1';
           if(RADDR <depth-1  ) then
             RADDR := RADDR + 1;
           else
             RADDR :=(RADDR +1) mod  depth;
             RADDR_wrap :=1 - RADDR_wrap;
           end if;
            do_par  := DO8_zd XOR DO7_zd XOR DO6_zd XOR DO5_zd XOR DO4_zd XOR DO3_zd XOR
                       DO2_zd XOR DO1_zd XOR DO0_zd;
            par_f <= do_par;
            if (do_par = 'X') then
             RPE_zd := 'X';
            elsif (do_par /= PARODD_delayed) then
             RPE_zd  :=  '1';
            else
             RPE_zd  :=  '0';
            end if;
         end if;
     when others =>
       if (TO_X01(RBint_previous) /= 'X') then
        assert false
        report ": RDB or RBLKB unknown"
        severity Error;
        end if;
           DO0_zd  := 'X';
           DO1_zd  := 'X';
           DO2_zd  := 'X';
           DO3_zd  := 'X';
           DO4_zd  := 'X';
           DO5_zd  := 'X';
           DO6_zd  := 'X';
           DO7_zd  := 'X';
           DO8_zd  := 'X';
     end case;
  elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='0') AND (TO_X01(RESET_delayed) = '1') AND (TO_X01(READ_AT_PREV_EDGE) = '1')) then
   READ_AT_PREV_EDGE <='0';
   if(RADDR = WADDR ) then
    if(RADDR_wrap = WADDR_wrap) then
       EMPTY_tmp := '1';
       FULL_tmp  := '0';
    end if;
   end if;
   if(RADDR /= WADDR ) then
    FULL_tmp  := '0';
   end if;
    if(WADDR_wrap = RADDR_wrap ) then
     if((WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((WADDR - RADDR) >= thresh  ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    else 
     if((depth + WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((depth + WADDR - RADDR) >= thresh ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    end if;
 else 
    null;
 end if;

   -- Mimic odd silicon flag behavior coming out of RESET with WB low
   
   if ( hold_full_low = 1 ) then
     FULL_zd := '0';
   else
     FULL_zd := FULL_tmp;
   end if;

   if ( hold_empty_low = 1 ) then
     EMPTY_zd := '0';
   elsif ( hold_empty_high = 1 ) then
     EMPTY_zd := '1';
   else
     EMPTY_zd := EMPTY_tmp;
   end if;

   if ( hold_eqth_high = 1 ) then
     EQTH_zd := '1';
   elsif ( hold_eqth_low = 1 ) then
     EQTH_zd := '0';
   else
     EQTH_zd := EQTH_tmp;
   end if;

   -- If LEVEL greater than DEPTH then GEQTH mimics FULL
   
   if ( hold_geqth_high = 1 ) then
     GEQTH_zd := '1';
   elsif ( hold_geqth_low = 1 ) then
     GEQTH_zd := '0';
   else
     if ( thresh > depth ) then
       GEQTH_zd := FULL_zd;
     else
       GEQTH_zd := GEQTH_tmp;
     end if;
   end if;


  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       WCLKS_previous  := WCLKS_ipd;
       RCLKS_previous   := RCLKS_ipd;
       RBint_previous   := RBint_delayed;
       RBint_delayed    := RBint;
       WBint_previous   := WBint_delayed;
       WBint_delayed    := WBint;
       DI0_delayed      := DI0_ipd;
       DI1_delayed      := DI1_ipd;
       DI2_delayed      := DI2_ipd;
       DI3_delayed      := DI3_ipd;
       DI4_delayed      := DI4_ipd;
       DI5_delayed      := DI5_ipd;
       DI6_delayed      := DI6_ipd;
       DI7_delayed      := DI7_ipd;
       DI8_delayed      := DI8_ipd;
       LGDEP0_previous  := LGDEP0_delayed;
       LGDEP0_delayed   := LGDEP0_ipd;
       LGDEP1_previous  := LGDEP1_delayed;
       LGDEP1_delayed   := LGDEP1_ipd;
       LGDEP2_previous  := LGDEP2_delayed;
       LGDEP2_delayed   := LGDEP2_ipd;
       LEVEL0_previous  := LEVEL0_delayed;
       LEVEL0_delayed   := LEVEL0_ipd;
       LEVEL1_previous  := LEVEL1_delayed;
       LEVEL1_delayed   := LEVEL1_ipd;
       LEVEL2_previous  := LEVEL2_delayed;
       LEVEL2_delayed   := LEVEL2_ipd;
       LEVEL3_previous  := LEVEL3_delayed;
       LEVEL3_delayed   := LEVEL3_ipd;
       LEVEL4_previous  := LEVEL4_delayed;
       LEVEL4_delayed   := LEVEL4_ipd;
       LEVEL5_previous  := LEVEL5_delayed;
       LEVEL5_delayed   := LEVEL5_ipd;
       LEVEL6_previous  := LEVEL6_delayed;
       LEVEL6_delayed   := LEVEL6_ipd;
       LEVEL7_previous  := LEVEL7_delayed;
       LEVEL7_delayed   := LEVEL7_ipd;
       PARODD_previous  := PARODD_delayed; 
       PARODD_delayed   := PARODD_ipd;
       RESET_previous   := RESET_delayed; 
       RESET_delayed    := RESET_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
             OutSignal     => DOS,
             GlitchData    => DOS_GlitchData,
             OutSignalName => "DOS",
             OutTemp       => DOS_zd,

             Paths =>   (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO0), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO1), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO2), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO3), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO4), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO5), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO6), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO7), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO8), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => FULL,
           GlitchData    => FULL_GlitchData,
           OutSignalName => "FULL",
           OutTemp       => FULL_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_FULL), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_FULL), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_FULL), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EMPTY,
           GlitchData    => EMPTY_GlitchData,
           OutSignalName => "EMPTY",
           OutTemp       => EMPTY_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EMPTY), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_EMPTY), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EMPTY), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EQTH,
           GlitchData    => EQTH_GlitchData,
           OutSignalName => "EQTH",
           OutTemp       => EQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EQTH), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_EQTH), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => GEQTH,
           GlitchData    => GEQTH_GlitchData,
           OutSignalName => "GEQTH",
           OutTemp       => GEQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_GEQTH), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_GEQTH), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_GEQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );


   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

LIBRARY a500k;
USE a500k.all;

entity FIFO256x9SSR is 
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_RPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_PARODD_WPE		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_WCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_WCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;

        -- WCLK falling edge setup to RESET rising edge 
 	trecovery_RESET_WCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_WCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- WCLK rising  edge hold to RESET rising edge 
	thold_RESET_WCLKS_posedge_posedge             : VitalDelayType := 0.00 ns;
	thold_RESET_WCLKS_posedge_negedge             : VitalDelayType := 0.00 ns;
	tpw_WCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        WPE    :  OUT STD_LOGIC := 'X';
        RPE    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        WCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');


ATTRIBUTE VITAL_LEVEL0 OF FIFO256x9SSR : entity IS True ;
END FIFO256x9SSR;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of FIFO256x9SSR is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal LGDEP0_ipd : std_ulogic := 'X';
   signal LGDEP1_ipd : std_ulogic := 'X';
   signal LGDEP2_ipd : std_ulogic := 'X';
   signal LEVEL0_ipd : std_ulogic := 'X';
   signal LEVEL1_ipd : std_ulogic := 'X';
   signal LEVEL2_ipd : std_ulogic := 'X';
   signal LEVEL3_ipd : std_ulogic := 'X';
   signal LEVEL4_ipd : std_ulogic := 'X';
   signal LEVEL5_ipd : std_ulogic := 'X';
   signal LEVEL6_ipd : std_ulogic := 'X';
   signal LEVEL7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal RESET_ipd  : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal WCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

   -- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic := 'X';
   signal par_f2     : std_logic := 'X';

   signal WRITE_AT_PREV_EDGE : std_logic := '0';
   signal READ_AT_PREV_EDGE  : std_logic := '0';

   begin  --  VITAL_ACT

   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (LGDEP0_ipd, LGDEP0, VitalExtendToFillDelay(tipd_LGDEP0));
   VitalWireDelay (LGDEP1_ipd, LGDEP1, VitalExtendToFillDelay(tipd_LGDEP1));
   VitalWireDelay (LGDEP2_ipd, LGDEP2, VitalExtendToFillDelay(tipd_LGDEP2));
   VitalWireDelay (LEVEL0_ipd, LEVEL0, VitalExtendToFillDelay(tipd_LEVEL0));
   VitalWireDelay (LEVEL1_ipd, LEVEL1, VitalExtendToFillDelay(tipd_LEVEL1));
   VitalWireDelay (LEVEL2_ipd, LEVEL2, VitalExtendToFillDelay(tipd_LEVEL2));
   VitalWireDelay (LEVEL3_ipd, LEVEL3, VitalExtendToFillDelay(tipd_LEVEL3));
   VitalWireDelay (LEVEL4_ipd, LEVEL4, VitalExtendToFillDelay(tipd_LEVEL4));
   VitalWireDelay (LEVEL5_ipd, LEVEL5, VitalExtendToFillDelay(tipd_LEVEL5));
   VitalWireDelay (LEVEL6_ipd, LEVEL6, VitalExtendToFillDelay(tipd_LEVEL6));
   VitalWireDelay (LEVEL7_ipd, LEVEL7, VitalExtendToFillDelay(tipd_LEVEL7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RESET_ipd, RESET, VitalExtendToFillDelay(tipd_RESET));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (WCLKS_ipd, WCLKS, VitalExtendToFillDelay(tipd_WCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

   ---------------------------------------------------------------
   --                  Behavior Section                         --
   ---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);

    VITALBehavior : process (
                          LEVEL0_ipd, LEVEL1_ipd, LEVEL2_ipd, LEVEL3_ipd, LEVEL4_ipd, LEVEL5_ipd, LEVEL6_ipd, LEVEL7_ipd, 
                          LGDEP0_ipd, LGDEP1_ipd, LGDEP2_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd, RESET_ipd
                          )

     -- some internal veriable declaration
     variable RAM_di_int   : std_logic_vector(8 downto 0);
     variable memory_array : MEM_TYPE  := (others =>(others => 'X'));
     variable do_par       : std_logic := 'X';
     variable tmp_par      : std_logic := 'X';
     variable tmp_par2     : std_logic := 'X';
     variable wpe_var      : std_logic := 'X';
     variable temp         : integer   := 0;
     variable thresh       : integer   := 0;
     variable depth        : integer   := 0;
     variable WADDR        : integer   := 0;
     variable WADDR_wrap   : integer   := 0;
     variable RADDR        : integer   := 0;
     variable RADDR_wrap   : integer   := 0;

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     --  Read Timing Check Results
     variable PeriodData_RESET           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET                : X01                 := '0';
     variable Tviol_PARODD_RCLKS_posedge : X01                 := '0';
     variable TmDt_PARODD_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_RCLKS_posedge  : X01                 := '0';
     variable Tmkr_RESET_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable Tviol_DI0_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI0_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI1_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI2_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI3_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI4_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI5_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI6_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI7_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI8_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_PARODD_WCLKS_posedge : X01                 := '0';
     variable TmDt_PARODD_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_WCLKS_posedge    : X01                 := '0';
     variable TmDt_WRB_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_WCLKS_posedge  : X01                 := '0';
     variable TmDt_WBLKB_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_WCLKS_posedge  : X01                 := '0';
     variable Tmkr_RESET_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WCLKS                : X01                 := '0';

     -- functional Results


     variable DO0_zd   : std_ulogic;
     variable DO1_zd   : std_ulogic;
     variable DO2_zd   : std_ulogic;
     variable DO3_zd   : std_ulogic;
     variable DO4_zd   : std_ulogic;
     variable DO5_zd   : std_ulogic;
     variable DO6_zd   : std_ulogic;
     variable DO7_zd   : std_ulogic;
     variable DO8_zd   : std_ulogic;
     variable RPE_zd   : std_ulogic;
     variable WPE_zd   : std_ulogic;
     variable DOS_zd   : std_ulogic;
     variable FULL_zd  : std_ulogic;
     variable EMPTY_zd : std_ulogic;
     variable EQTH_zd  : std_ulogic;
     variable GEQTH_zd : std_ulogic;
     variable FULL_tmp  : std_ulogic;
     variable EMPTY_tmp : std_ulogic;
     variable EQTH_tmp  : std_ulogic;
     variable GEQTH_tmp : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData   : VitalGlitchDataType;
     variable DO1_GlitchData   : VitalGlitchDataType;
     variable DO2_GlitchData   : VitalGlitchDataType;
     variable DO3_GlitchData   : VitalGlitchDataType;
     variable DO4_GlitchData   : VitalGlitchDataType;
     variable DO5_GlitchData   : VitalGlitchDataType;
     variable DO6_GlitchData   : VitalGlitchDataType;
     variable DO7_GlitchData   : VitalGlitchDataType;
     variable DO8_GlitchData   : VitalGlitchDataType;
     variable RPE_GlitchData   : VitalGlitchDataType;
     variable WPE_GlitchData   : VitalGlitchDataType;
     variable DOS_GlitchData   : VitalGlitchDataType;
     variable FULL_GlitchData  : VitalGlitchDataType;
     variable EMPTY_GlitchData : VitalGlitchDataType;
     variable EQTH_GlitchData  : VitalGlitchDataType;
     variable GEQTH_GlitchData : VitalGlitchDataType;

     -- last value variables
     variable WCLKS_previous   : std_ulogic := 'X';
     variable RCLKS_previous   : std_ulogic := 'X';
     variable RBint_delayed    : std_ulogic := 'X';
     variable RBint_previous   : std_ulogic := 'X';
     variable WBint_delayed    : std_ulogic := 'X';
     variable WBint_previous   : std_ulogic := 'X';
     variable DIS_previous     : std_ulogic := 'X';
     variable RESET_previous   : std_ulogic := 'X';
     variable RESET_delayed    : std_ulogic := 'X';
     variable PARODD_previous  : std_ulogic := 'X';
     variable PARODD_delayed   : std_ulogic := 'X';
     variable DI0_delayed      : std_ulogic := 'X';
     variable DI1_delayed      : std_ulogic := 'X';
     variable DI2_delayed      : std_ulogic := 'X';
     variable DI3_delayed      : std_ulogic := 'X';
     variable DI4_delayed      : std_ulogic := 'X';
     variable DI5_delayed      : std_ulogic := 'X';
     variable DI6_delayed      : std_ulogic := 'X';
     variable DI7_delayed      : std_ulogic := 'X';
     variable DI8_delayed      : std_ulogic := 'X';
     variable DI0_previous     : std_ulogic := 'X';
     variable DI1_previous     : std_ulogic := 'X';
     variable DI2_previous     : std_ulogic := 'X';
     variable DI3_previous     : std_ulogic := 'X';
     variable DI4_previous     : std_ulogic := 'X';
     variable DI5_previous     : std_ulogic := 'X';
     variable DI6_previous     : std_ulogic := 'X';
     variable DI7_previous     : std_ulogic := 'X';
     variable DI8_previous     : std_ulogic := 'X';
     variable LGDEP0_delayed   : std_ulogic := 'X';
     variable LGDEP1_delayed   : std_ulogic := 'X';
     variable LGDEP2_delayed   : std_ulogic := 'X';
     variable LGDEP0_previous  : std_ulogic := 'X';
     variable LGDEP1_previous  : std_ulogic := 'X';
     variable LGDEP2_previous  : std_ulogic := 'X';
     variable LEVEL0_delayed   : std_ulogic := 'X';
     variable LEVEL1_delayed   : std_ulogic := 'X';
     variable LEVEL2_delayed   : std_ulogic := 'X';
     variable LEVEL3_delayed   : std_ulogic := 'X';
     variable LEVEL4_delayed   : std_ulogic := 'X';
     variable LEVEL5_delayed   : std_ulogic := 'X';
     variable LEVEL6_delayed   : std_ulogic := 'X';
     variable LEVEL7_delayed   : std_ulogic := 'X';
     variable LEVEL0_previous  : std_ulogic := 'X';
     variable LEVEL1_previous  : std_ulogic := 'X';
     variable LEVEL2_previous  : std_ulogic := 'X';
     variable LEVEL3_previous  : std_ulogic := 'X';
     variable LEVEL4_previous  : std_ulogic := 'X';
     variable LEVEL5_previous  : std_ulogic := 'X';
     variable LEVEL6_previous  : std_ulogic := 'X';
     variable LEVEL7_previous  : std_ulogic := 'X';

     --  Pipelined temporary results
     variable RPE_stg1         : std_ulogic := 'X';
     variable DO0_stg1         : std_ulogic := 'X';
     variable DO1_stg1         : std_ulogic := 'X';
     variable DO2_stg1         : std_ulogic := 'X';
     variable DO3_stg1         : std_ulogic := 'X';
     variable DO4_stg1         : std_ulogic := 'X';
     variable DO5_stg1         : std_ulogic := 'X';
     variable DO6_stg1         : std_ulogic := 'X';
     variable DO7_stg1         : std_ulogic := 'X';
     variable DO8_stg1         : std_ulogic := 'X';

     -- Special variables to control flags
     variable hold_empty_low   : integer := 0;
     variable hold_eqth_high   : integer := 0;
     variable hold_geqth_high  : integer := 0;
     variable hold_full_low    : integer := 0;
     variable hold_empty_high  : integer := 0;
     variable hold_eqth_low    : integer := 0;
     variable hold_geqth_low   : integer := 0;

     variable WCLKS_re         : Time;
     variable WCLKS_fe         : Time;
     variable WCLKS_fe_prev    : Time;
     variable WB_re            : Time;
     variable RESET_re         : Time;

 begin -- process VITALBehavior

 if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

   -- recovery / removal check for RCLKS to RESET signal ;
       VitalRecoveryRemovalCheck ( Tviol_RESET_RCLKS_posedge,
                             Tmkr_RESET_RCLKS_posedge,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             trecovery_RESET_RCLKS_posedge_negedge,
                             thold_RESET_RCLKS_posedge_posedge,
                             TRUE,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'), 
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             TRUE,
                             TRUE,
                             WARNING
                             );

   -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             ((TO_X01(RBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             ((TO_X01(RDB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_PARODD_RCLKS_posedge,
                             TmDt_PARODD_RCLKS_posedge,
                             PARODD_ipd, "PARODD",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_PARODD_RCLKS_posedge_posedge,
                             tsetup_PARODD_RCLKS_negedge_posedge,
                             thold_PARODD_RCLKS_posedge_posedge,
                             thold_PARODD_RCLKS_negedge_posedge,
                             (TO_X01(RESET_ipd) = '1'),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (TO_X01(RDB) = '0') AND (TO_X01(RBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9SSR",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RESET,
                              PeriodData_RESET,
                              RESET_ipd, "RESET",
                              0.0 ns,
                              tpw_RESET_negedge,
                              0.0 ns,
                              tpw_RESET_negedge,
                              True,
                              InstancePath & "/FIFO256x9SSR",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       -- recovery / removal check for WCLKS to RESET signal ;
       VitalRecoveryRemovalCheck ( Tviol_RESET_WCLKS_posedge,
                             Tmkr_RESET_WCLKS_posedge,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns,
                             trecovery_RESET_WCLKS_posedge_negedge,
                             thold_RESET_WCLKS_posedge_posedge,
                             TRUE,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'), 
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             TRUE,
                             TRUE,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_posedge_posedge,
                             tsetup_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_posedge_posedge,
                             tsetup_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_posedge_posedge,
                             tsetup_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_posedge_posedge,
                             tsetup_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_posedge_posedge,
                             tsetup_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_posedge_posedge,
                             tsetup_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_posedge_posedge,
                             tsetup_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_posedge_posedge,
                             tsetup_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_posedge_posedge,
                             tsetup_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

   -- setup hold WEN, WBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_posedge_posedge,
                             tsetup_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_PARODD_WCLKS_posedge,
                             TmDt_PARODD_WCLKS_posedge,
                             PARODD_ipd, "PARODD",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_PARODD_WCLKS_posedge_posedge,
                             tsetup_PARODD_WCLKS_negedge_posedge,
                             thold_PARODD_WCLKS_posedge_posedge,
                             thold_PARODD_WCLKS_negedge_posedge,
                             ((TO_X01(RBint) = '0') AND (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/FIFO256x9SSR",
                             True,
                             True,
                             WARNING
                             );

  --   Period of WCLK
      VitalPeriodPulseCheck ( Pviol_WCLKS,
                              PeriodData_WCLKS,
                              WCLKS_ipd, "WCLKS",
                              0.0 ns,
                              tperiod_WCLKS,
                              tpw_WCLKS_posedge,
                              tpw_WCLKS_negedge,
                              (TO_X01(WRB) = '0') AND (TO_X01(WBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9SSR",
                              True,
                              True,
                              WARNING
                              );
 end if;

   ------------------------------------------------------------
   --               FIFO RESET                               --
   ------------------------------------------------------------

   if ( RESET_ipd'event and RESET_ipd = '0' ) then
       WADDR      := 0;
       RADDR      := 0;
       WADDR_wrap := 0;
       RADDR_wrap := 0;
       FULL_tmp   := '0';
       EMPTY_tmp  := '1';
       EQTH_tmp   := '0';
       GEQTH_tmp  := '0';
       WRITE_AT_PREV_EDGE <='0';
       READ_AT_PREV_EDGE <='0';
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
       hold_full_low   := 0;
       hold_empty_high := 0;
       hold_eqth_low   := 0;
       hold_geqth_low  := 0;
   end if;

   if ( WCLKS_ipd'event and WCLKS_ipd = '1' ) then
     WCLKS_re := now;
   end if;
      
   if ( WBint'event and WBint = '1' ) then
     WB_re := now;
   end if;
      
   if ( RESET_ipd'event and RESET_ipd = '1' ) then
     RESET_re := now;
     if ( TO_X01 ( WCLKS_ipd ) = '1' ) then
       if ( WCLKS_re = WB_re ) then
         hold_full_low   := 1; -- until next reset
         hold_empty_high := 1;
         hold_eqth_low   := 1;
         hold_geqth_low  := 1;
       elsif ( TO_X01 ( WBint ) = '0' ) then
         EMPTY_zd        := '0';
         EQTH_zd         := '1';
         GEQTH_zd        := '1';
         hold_empty_low  := 1; -- until next WCLKS falling edge
         hold_eqth_high  := 1;
         hold_geqth_high := 1;
       elsif ( WCLKS_re < WB_re ) then
         EMPTY_zd        := '0';
         EQTH_zd         := '1';
         GEQTH_zd        := '1';
         hold_empty_low  := 1; -- until next WCLKS falling edge
         hold_eqth_high  := 1;
         hold_geqth_high := 1;
       elsif ( WB_re < WCLKS_re ) then
         hold_empty_low  := 0; -- expected behavior
         hold_eqth_high  := 0;
         hold_geqth_high := 0;
         hold_full_low   := 0;
         hold_empty_high := 0;
         hold_eqth_low   := 0;
         hold_geqth_low  := 0;
       end if;
     else
       hold_empty_low  := 0; -- expected behavior
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
       hold_full_low   := 0;
       hold_empty_high := 0;
       hold_eqth_low   := 0;
       hold_geqth_low  := 0;
     end if;
   end if;

   if ( WCLKS_ipd'event and WCLKS_ipd = '0' ) then
     WCLKS_fe_prev := WCLKS_fe;
     WCLKS_fe := now;
     if (( TO_X01 ( RESET_ipd ) = '1' ) and ( WCLKS_fe_prev < RESET_re )) then
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
     end if;
   end if;

   ------------------------------------------------------------
   -- WPE output                                              -
   ------------------------------------------------------------

   if ( PARODD_ipd'EVENT ) then
     RPE_zd := not RPE_zd;
     WPE_zd := not WPE_zd;
     RPE_stg1 := not RPE_stg1;
   end if;

   ------------------------------------------------------------
   --         WPE generating block                            -
   ------------------------------------------------------------

    if (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
        tmp_par := DI7_delayed XOR DI6_delayed XOR DI5_delayed XOR DI4_delayed XOR DI3_delayed XOR DI2_delayed XOR DI1_delayed XOR DI0_delayed;
        par_f    <= tmp_par ;
        tmp_par2 := (tmp_par xor DI8_delayed);
        par_f2   <= tmp_par2;

      if (( TO_X01 ( PARODD_ipd ) = 'X' ) or 
          ( TO_X01 ( DI8_ipd )    = 'X' ) or
          ( TO_X01 ( DI7_ipd )    = 'X' ) or
          ( TO_X01 ( DI6_ipd )    = 'X' ) or
          ( TO_X01 ( DI5_ipd )    = 'X' ) or
          ( TO_X01 ( DI4_ipd )    = 'X' ) or
          ( TO_X01 ( DI3_ipd )    = 'X' ) or
          ( TO_X01 ( DI2_ipd )    = 'X' ) or
          ( TO_X01 ( DI1_ipd )    = 'X' ) or
          ( TO_X01 ( DI0_ipd )    = 'X' )
         ) then
        wpe_var  :=  'X';
      else
        if ( tmp_par2 /= PARODD_ipd ) then
          wpe_var  :=  '1';
        else
          wpe_var  :=  '0';
        end if;
      end if;

        RAM_di_int(8) := DI8_delayed;
        WPE_zd := wpe_var;
    end if;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

   if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
   end if; 

   -----------------------------------------------------------
   --    calculate the depth and levels                     --
   -----------------------------------------------------------

    temp :=((INT(LGDEP2_delayed)*4) + (INT(LGDEP1_delayed)*2) + 
           (INT(LGDEP0_delayed)*1));

    case temp is 
         when 0 => depth := 2;
         when 1 => depth := 4;
         when 2 => depth := 8;
         when 3 => depth := 16;
         when 4 => depth := 32;
         when 5 => depth := 64;
         when 6 => depth := 128;
         when 7 => depth := 256;
         when others => depth := 0;
    end case;

    -- thresh value

    thresh := (INT(LEVEL7_delayed)*128) + (INT(LEVEL6_delayed)*64) + 
               (INT(LEVEL5_delayed)*32) + (INT(LEVEL4_delayed)*16) + 
               (INT(LEVEL3_delayed)*8) + (INT(LEVEL2_delayed)*4) + 
               (INT(LEVEL1_delayed)*2) + (INT(LEVEL0_delayed)*1); 

    if ( thresh = 0 or thresh = 255 ) then
      assert false
        report " Illegal level configuration, LEVEL cannot be 0 or 255 "
        severity failure;
    end if;

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

   if(TO_X01(WCLKS_ipd)='X') then
    if(RESET_delayed = '1') then
     if (WBint_delayed = '0') then
      if (TO_X01(WCLKS_previous) /= 'X') then
        assert false
        report ": WCLK unknown"
        severity Error;
      end if;
     end if;
    end if;
   elsif (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') AND (TO_X01(RESET_ipd) = '1')then
     WRITE_AT_PREV_EDGE <='0';
     case (TO_X01(WBint_delayed)) is 
      when '1' =>
                null;
      when '0' => 
         if(FULL_zd = '0') then 
         RAM_di_int(7 downto 0) := DI7_delayed & DI6_delayed & DI5_delayed & 
                                    DI4_delayed & DI3_delayed & DI2_delayed & 
                                    DI1_delayed & DI0_delayed;
         memory_array(WADDR) := RAM_di_int;
         WRITE_AT_PREV_EDGE <='1';
         if(WADDR <depth-1  ) then
           WADDR := WADDR + 1;
         elsif( WADDR  = depth-1) then
           WADDR := 0;
           WADDR_wrap := 1 - WADDR_wrap;
         end if;
        end if;
       when others => 
        if (TO_X01(WBint_previous) /= 'X') then
          assert false
          report ": WBLKB or WRB unknown"
          severity Error;
          end if;
        end case;
     elsif(WCLKS_ipd'EVENT AND WCLKS_ipd = '0')  AND (TO_X01(RESET_delayed) = '1') AND (TO_X01(WRITE_AT_PREV_EDGE) = '1')then
        WRITE_AT_PREV_EDGE <='0';
        if(WADDR   = RADDR ) then
         if(RADDR_wrap /= WADDR_wrap) then
          FULL_tmp := '1';
          EMPTY_tmp :='0';
         end if;
        end if;
        if(WADDR   /= RADDR ) then
          EMPTY_tmp := '0';
        end if;
          if(RADDR_wrap = WADDR_wrap) then
            if(WADDR - RADDR = thresh ) then
               EQTH_tmp := '1';
            else 
               EQTH_tmp := '0';
            end if;
            if(WADDR - RADDR >= thresh ) then
                GEQTH_tmp := '1';
            else 
                GEQTH_tmp := '0';
            end if;
          else 
           if((depth -RADDR + WADDR) = thresh ) then
               EQTH_tmp := '1';
            else 
               EQTH_tmp := '0';
            end if;
            if((depth -RADDR + WADDR) >= thresh ) then
                GEQTH_tmp := '1';
            else 
                GEQTH_tmp := '0';
            end if;
           end if; 
      else
       null;
    end if;


  --------------------------------------------------------------------
  --          FIFO READ SECTION........                             --
  --------------------------------------------------------------------

  if (TO_X01(RCLKS_ipd)='X') then
    if(RESET_ipd /= '0') then
    if(TO_X01(RBint_delayed) /= '1') then
      if(TO_X01(RCLKS_previous) /= 'X') then
        assert false
        report ": RCLK unknown"
        severity Error;
        DO0_zd  := 'X';
        DO1_zd  := 'X';
        DO2_zd  := 'X';
        DO3_zd  := 'X';
        DO4_zd  := 'X';
        DO5_zd  := 'X';
        DO6_zd  := 'X';
        DO7_zd  := 'X';
        DO8_zd  := 'X';
      end if;
     end if;
    end if;
   elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='1') AND (TO_X01(RESET_delayed) = '1')) then
     DO0_zd := DO0_stg1;
     DO1_zd := DO1_stg1;
     DO2_zd := DO2_stg1;
     DO3_zd := DO3_stg1;
     DO4_zd := DO4_stg1;
     DO5_zd := DO5_stg1;
     DO6_zd := DO6_stg1;
     DO7_zd := DO7_stg1;
     DO8_zd := DO8_stg1;
     RPE_zd := RPE_stg1;
     READ_AT_PREV_EDGE <='0';
     case (TO_X01(RBint_delayed)) is
        when '1' =>
                null;
        when '0' =>
         if(TO_X01(EMPTY_zd) /= '1') then 
           DO0_stg1  := memory_array(RADDR)(0);
           DO1_stg1  := memory_array(RADDR)(1);
           DO2_stg1  := memory_array(RADDR)(2);
           DO3_stg1  := memory_array(RADDR)(3);
           DO4_stg1  := memory_array(RADDR)(4);
           DO5_stg1  := memory_array(RADDR)(5);
           DO6_stg1  := memory_array(RADDR)(6);
           DO7_stg1  := memory_array(RADDR)(7);
           DO8_stg1  := memory_array(RADDR)(8);
           READ_AT_PREV_EDGE <='1';
           if(RADDR <depth-1  ) then
             RADDR := RADDR + 1;
           else
             RADDR :=(RADDR +1) mod  depth;
             RADDR_wrap :=1 - RADDR_wrap;
           end if;
      do_par  := DO8_stg1 XOR DO7_stg1 XOR DO6_stg1 XOR DO5_stg1 XOR DO4_stg1 XOR DO3_stg1 XOR
                 DO2_stg1 XOR DO1_stg1 XOR DO0_stg1;
            par_f <= do_par;
            if (do_par = 'X') then
             RPE_stg1 := 'X';
            elsif (do_par /= PARODD_delayed) then
             RPE_stg1  :=  '1';
            else
             RPE_stg1  :=  '0';
            end if;
         end if;
     when others =>
       if (TO_X01(RBint_previous) /= 'X') then
        assert false
        report ": RDB or RBLKB unknown"
        severity Error;
        end if;
           DO0_stg1  := 'X';
           DO1_stg1  := 'X';
           DO2_stg1  := 'X';
           DO3_stg1  := 'X';
           DO4_stg1  := 'X';
           DO5_stg1  := 'X';
           DO6_stg1  := 'X';
           DO7_stg1  := 'X';
           DO8_stg1  := 'X';
     end case;
  elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='0') AND (TO_X01(RESET_delayed) = '1') AND (TO_X01(READ_AT_PREV_EDGE) = '1')) then
   READ_AT_PREV_EDGE <='0';
   if(RADDR = WADDR ) then
    if(RADDR_wrap = WADDR_wrap) then
       EMPTY_tmp := '1';
       FULL_tmp  := '0';
    end if;
   end if;
   if(RADDR /= WADDR ) then
    FULL_tmp  := '0';
   end if;
    if(WADDR_wrap = RADDR_wrap ) then
     if((WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((WADDR - RADDR) >= thresh  ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    else 
     if((depth + WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((depth + WADDR - RADDR) >= thresh ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    end if;
 else 
    null;
 end if;

   -- Mimic odd silicon flag behavior coming out of RESET with WB low
   
   if ( hold_full_low = 1 ) then
     FULL_zd := '0';
   else
     FULL_zd := FULL_tmp;
   end if;

   if ( hold_empty_low = 1 ) then
     EMPTY_zd := '0';
   elsif ( hold_empty_high = 1 ) then
     EMPTY_zd := '1';
   else
     EMPTY_zd := EMPTY_tmp;
   end if;

   if ( hold_eqth_high = 1 ) then
     EQTH_zd := '1';
   elsif ( hold_eqth_low = 1 ) then
     EQTH_zd := '0';
   else
     EQTH_zd := EQTH_tmp;
   end if;

   -- If LEVEL greater than DEPTH then GEQTH mimics FULL
   
   if ( hold_geqth_high = 1 ) then
     GEQTH_zd := '1';
   elsif ( hold_geqth_low = 1 ) then
     GEQTH_zd := '0';
   else
     if ( thresh > depth ) then
       GEQTH_zd := FULL_zd;
     else
       GEQTH_zd := GEQTH_tmp;
     end if;
   end if;


  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       WCLKS_previous  := WCLKS_ipd;
       RCLKS_previous   := RCLKS_ipd;
       RBint_previous   := RBint_delayed;
       RBint_delayed    := RBint;
       WBint_previous   := WBint_delayed;
       WBint_delayed    := WBint;
       DI0_delayed      := DI0_ipd;
       DI1_delayed      := DI1_ipd;
       DI2_delayed      := DI2_ipd;
       DI3_delayed      := DI3_ipd;
       DI4_delayed      := DI4_ipd;
       DI5_delayed      := DI5_ipd;
       DI6_delayed      := DI6_ipd;
       DI7_delayed      := DI7_ipd;
       DI8_delayed      := DI8_ipd;
       LGDEP0_previous  := LGDEP0_delayed;
       LGDEP0_delayed   := LGDEP0_ipd;
       LGDEP1_previous  := LGDEP1_delayed;
       LGDEP1_delayed   := LGDEP1_ipd;
       LGDEP2_previous  := LGDEP2_delayed;
       LGDEP2_delayed   := LGDEP2_ipd;
       LEVEL0_previous  := LEVEL0_delayed;
       LEVEL0_delayed   := LEVEL0_ipd;
       LEVEL1_previous  := LEVEL1_delayed;
       LEVEL1_delayed   := LEVEL1_ipd;
       LEVEL2_previous  := LEVEL2_delayed;
       LEVEL2_delayed   := LEVEL2_ipd;
       LEVEL3_previous  := LEVEL3_delayed;
       LEVEL3_delayed   := LEVEL3_ipd;
       LEVEL4_previous  := LEVEL4_delayed;
       LEVEL4_delayed   := LEVEL4_ipd;
       LEVEL5_previous  := LEVEL5_delayed;
       LEVEL5_delayed   := LEVEL5_ipd;
       LEVEL6_previous  := LEVEL6_delayed;
       LEVEL6_delayed   := LEVEL6_ipd;
       LEVEL7_previous  := LEVEL7_delayed;
       LEVEL7_delayed   := LEVEL7_ipd;
       PARODD_previous  := PARODD_delayed; 
       PARODD_delayed   := PARODD_ipd;
       RESET_previous   := RESET_delayed; 
       RESET_delayed    := RESET_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
             OutSignal     => DOS,
             GlitchData    => DOS_GlitchData,
             OutSignalName => "DOS",
             OutTemp       => DOS_zd,

             Paths =>   (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
           OutSignal     => WPE,
           GlitchData    => WPE_GlitchData,
           OutSignalName => "WPE",
           OutTemp       => WPE_zd,
           Paths =>   (0  => (WCLKS_ipd'last_event,
                       VitalExtendToFillDelay(tpd_WCLKS_WPE), true),
                       1 => (PARODD_ipd'last_event,
                             VitalExtendToFillDelay(tpd_PARODD_WPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO0), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO1), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO2), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO3), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO4), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO5), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO6), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO7), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO8), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => RPE,
           GlitchData    => RPE_GlitchData,
           OutSignalName => "RPE",
           OutTemp       => RPE_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_RPE), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_RPE), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => FULL,
           GlitchData    => FULL_GlitchData,
           OutSignalName => "FULL",
           OutTemp       => FULL_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_FULL), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_FULL), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_FULL), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EMPTY,
           GlitchData    => EMPTY_GlitchData,
           OutSignalName => "EMPTY",
           OutTemp       => EMPTY_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EMPTY), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_EMPTY), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EMPTY), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EQTH,
           GlitchData    => EQTH_GlitchData,
           OutSignalName => "EQTH",
           OutTemp       => EQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EQTH), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_EQTH), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => GEQTH,
           GlitchData    => GEQTH_GlitchData,
           OutSignalName => "GEQTH",
           OutTemp       => GEQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_GEQTH), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_GEQTH), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_GEQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );


   end process VITALBehavior;

  end VITAL_ACT;


LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
USE ieee.std_logic_unsigned.all;
USE IEEE.VITAL_timing.all;
USE IEEE.VITAL_primitives.all;

LIBRARY a500k;
USE a500k.all;

entity FIFO256x9SSRP is 
   generic (
        Xon           : Boolean := False;
        MsgOn         : Boolean := True;
        TimingCheckOn : Boolean := True;
        InstancePath  : String  := "*";

 	tipd_LEVEL0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LEVEL7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_LGDEP2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RCLKS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WRB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RDB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_WBLKB		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DIS		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_PARODD		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_RESET		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI0		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI1		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI2		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI3		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI4		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI5		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI6		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI7		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tipd_DI8		: VitalDelayType01Z     := (0 ns, 0 ns, 0 ns, 0 ns, 0 ns, 0 ns);
 	tpd_DIS_DOS		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
	tpd_WCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RCLKS_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_FULL		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EMPTY		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_EQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_GEQTH		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO0		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO1		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO2		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO3		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO4		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO5		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO6		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO7		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);
 	tpd_RESET_DO8		: VitalDelayType01Z     := (0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns, 0.1 ns);

 	tsetup_RDB_RCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_RDB_RCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_RBLKB_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_RBLKB_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_RCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_RCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	thold_RDB_RCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_RDB_RCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_RBLKB_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RBLKB_RCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_RCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_RCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;

        -- RCLK falling edge setup to RESET rising edge 
	trecovery_RESET_RCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_RCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- RCLK rising  edge hold to RESET rising edge 
 	thold_RESET_RCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_RESET_RCLKS_posedge_negedge             : VitalDelayType := 0.000 ns;
	tpw_RCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_RCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_RCLKS                                 : VitalDelayType := 0.000 ns;

 	tpw_RESET_negedge                             : VitalDelayType := 0.000 ns;
 	tsetup_WRB_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_WRB_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_WBLKB_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
	tsetup_WBLKB_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
 	tsetup_PARODD_WCLKS_posedge_posedge           : VitalDelayType := 0.000 ns;
	tsetup_PARODD_WCLKS_negedge_posedge           : VitalDelayType := 0.000 ns;
 	tsetup_DI0_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI0_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI1_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI1_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI2_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI2_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI3_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI3_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI4_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI4_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI5_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI5_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI6_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI6_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI7_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI7_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	tsetup_DI8_WCLKS_posedge_posedge              : VitalDelayType := 0.000 ns;
	tsetup_DI8_WCLKS_negedge_posedge              : VitalDelayType := 0.000 ns;
 	thold_WRB_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_WRB_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_WBLKB_WCLKS_posedge_posedge             : VitalDelayType := 0.000 ns;
	thold_WBLKB_WCLKS_negedge_posedge             : VitalDelayType := 0.000 ns;
 	thold_PARODD_WCLKS_negedge_posedge            : VitalDelayType := 0.000 ns;
	thold_PARODD_WCLKS_posedge_posedge            : VitalDelayType := 0.000 ns;
 	thold_DI0_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI0_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI1_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI1_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI2_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI2_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI3_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI3_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI4_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI4_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI5_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI5_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI6_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI6_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI7_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI7_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;
 	thold_DI8_WCLKS_posedge_posedge               : VitalDelayType := 0.000 ns;
	thold_DI8_WCLKS_negedge_posedge               : VitalDelayType := 0.000 ns;

        -- WCLK falling edge setup to RESET rising edge 
 	trecovery_RESET_WCLKS_posedge_posedge            : VitalDelayType := 0.00 ns;
	trecovery_RESET_WCLKS_posedge_negedge            : VitalDelayType := 0.00 ns;

        -- WCLK rising  edge hold to RESET rising edge 
	thold_RESET_WCLKS_posedge_posedge             : VitalDelayType := 0.00 ns;
	thold_RESET_WCLKS_posedge_negedge             : VitalDelayType := 0.00 ns;
	tpw_WCLKS_posedge                             : VitalDelayType := 0.000 ns;
 	tpw_WCLKS_negedge                             : VitalDelayType := 0.000 ns;
 	tperiod_WCLKS                                 : VitalDelayType := 0.000 ns
 	);

   port (
        DO0    :  OUT STD_LOGIC := 'X';
        DO1    :  OUT STD_LOGIC := 'X';
        DO2    :  OUT STD_LOGIC := 'X';
        DO3    :  OUT STD_LOGIC := 'X';
        DO4    :  OUT STD_LOGIC := 'X';
        DO5    :  OUT STD_LOGIC := 'X';
        DO6    :  OUT STD_LOGIC := 'X';
        DO7    :  OUT STD_LOGIC := 'X';
        DO8    :  OUT STD_LOGIC := 'X';
        DOS    :  OUT STD_LOGIC := 'X';
        FULL   :  OUT STD_LOGIC := 'X';
        EMPTY  :  OUT STD_LOGIC := 'X';
        EQTH   :  OUT STD_LOGIC := 'X';
        GEQTH  :  OUT STD_LOGIC := 'X';

        LGDEP0 :  IN STD_LOGIC := 'X';
        LGDEP1 :  IN STD_LOGIC := 'X';
        LGDEP2 :  IN STD_LOGIC := 'X';
        LEVEL0 :  IN STD_LOGIC := 'X';
        LEVEL1 :  IN STD_LOGIC := 'X';
        LEVEL2 :  IN STD_LOGIC := 'X';
        LEVEL3 :  IN STD_LOGIC := 'X';
        LEVEL4 :  IN STD_LOGIC := 'X';
        LEVEL5 :  IN STD_LOGIC := 'X';
        LEVEL6 :  IN STD_LOGIC := 'X';
        LEVEL7 :  IN STD_LOGIC := 'X';
        DI0    :  IN STD_LOGIC := 'X';
        DI1    :  IN STD_LOGIC := 'X';
        DI2    :  IN STD_LOGIC := 'X';
        DI3    :  IN STD_LOGIC := 'X';
        DI4    :  IN STD_LOGIC := 'X';
        DI5    :  IN STD_LOGIC := 'X';
        DI6    :  IN STD_LOGIC := 'X';
        DI7    :  IN STD_LOGIC := 'X';
        DI8    :  IN STD_LOGIC := 'X';
        WRB    :  IN STD_LOGIC := 'X';
        RDB    :  IN STD_LOGIC := 'X';
        WBLKB  :  IN STD_LOGIC := 'X';
        RBLKB  :  IN STD_LOGIC := 'X';
        PARODD :  IN STD_LOGIC := 'X';
        RESET  :  IN STD_LOGIC := 'X';
        RCLKS  :  IN STD_LOGIC := 'X';
        WCLKS  :  IN STD_LOGIC := 'X';
        DIS    :  IN STD_LOGIC := 'X');


ATTRIBUTE VITAL_LEVEL0 OF FIFO256x9SSRP : entity IS True ;
END FIFO256x9SSRP;



------------------------------------------------------
--  ARCHITECTURE declaration
------------------------------------------------------

architecture VITAL_ACT of FIFO256x9SSRP is

   attribute VITAL_LEVEL1 of VITAL_ACT : architecture is FALSE;

   signal LGDEP0_ipd : std_ulogic := 'X';
   signal LGDEP1_ipd : std_ulogic := 'X';
   signal LGDEP2_ipd : std_ulogic := 'X';
   signal LEVEL0_ipd : std_ulogic := 'X';
   signal LEVEL1_ipd : std_ulogic := 'X';
   signal LEVEL2_ipd : std_ulogic := 'X';
   signal LEVEL3_ipd : std_ulogic := 'X';
   signal LEVEL4_ipd : std_ulogic := 'X';
   signal LEVEL5_ipd : std_ulogic := 'X';
   signal LEVEL6_ipd : std_ulogic := 'X';
   signal LEVEL7_ipd : std_ulogic := 'X';
   signal DI0_ipd    : std_ulogic := 'X';
   signal DI1_ipd    : std_ulogic := 'X';
   signal DI2_ipd    : std_ulogic := 'X';
   signal DI3_ipd    : std_ulogic := 'X';
   signal DI4_ipd    : std_ulogic := 'X';
   signal DI5_ipd    : std_ulogic := 'X';
   signal DI6_ipd    : std_ulogic := 'X';
   signal DI7_ipd    : std_ulogic := 'X';
   signal DI8_ipd    : std_ulogic := 'X';
   signal RESET_ipd  : std_ulogic := 'X';
   signal WRB_ipd    : std_ulogic := 'X';
   signal RDB_ipd    : std_ulogic := 'X';
   signal WBLKB_ipd  : std_ulogic := 'X';
   signal RBLKB_ipd  : std_ulogic := 'X';
   signal PARODD_ipd : std_ulogic := 'X';
   signal RCLKS_ipd  : std_ulogic := 'X';
   signal WCLKS_ipd  : std_ulogic := 'X';
   signal DIS_ipd    : std_ulogic := 'X';

   -- New internal signals required
   signal WBint      : std_ulogic := 'X';
   signal RBint      : std_ulogic := 'X';

   TYPE MEM_TYPE IS ARRAY (255 DOWNTO 0) OF STD_LOGIC_VECTOR (8 DOWNTO 0);

   signal par_f      : std_logic := 'X';
   signal par_f2     : std_logic := 'X';

   signal WRITE_AT_PREV_EDGE : std_logic := '0';
   signal READ_AT_PREV_EDGE  : std_logic := '0';

   begin  --  VITAL_ACT

   --------------------------------------------------------
   --  INPUT PATH DELAYS                                 --
   --------------------------------------------------------

   WIRE_DELAY: block
   begin --  block WIRE_DELAY

   VitalWireDelay (LGDEP0_ipd, LGDEP0, VitalExtendToFillDelay(tipd_LGDEP0));
   VitalWireDelay (LGDEP1_ipd, LGDEP1, VitalExtendToFillDelay(tipd_LGDEP1));
   VitalWireDelay (LGDEP2_ipd, LGDEP2, VitalExtendToFillDelay(tipd_LGDEP2));
   VitalWireDelay (LEVEL0_ipd, LEVEL0, VitalExtendToFillDelay(tipd_LEVEL0));
   VitalWireDelay (LEVEL1_ipd, LEVEL1, VitalExtendToFillDelay(tipd_LEVEL1));
   VitalWireDelay (LEVEL2_ipd, LEVEL2, VitalExtendToFillDelay(tipd_LEVEL2));
   VitalWireDelay (LEVEL3_ipd, LEVEL3, VitalExtendToFillDelay(tipd_LEVEL3));
   VitalWireDelay (LEVEL4_ipd, LEVEL4, VitalExtendToFillDelay(tipd_LEVEL4));
   VitalWireDelay (LEVEL5_ipd, LEVEL5, VitalExtendToFillDelay(tipd_LEVEL5));
   VitalWireDelay (LEVEL6_ipd, LEVEL6, VitalExtendToFillDelay(tipd_LEVEL6));
   VitalWireDelay (LEVEL7_ipd, LEVEL7, VitalExtendToFillDelay(tipd_LEVEL7));
   VitalWireDelay (DI0_ipd, DI0, VitalExtendToFillDelay(tipd_DI0));
   VitalWireDelay (DI1_ipd, DI1, VitalExtendToFillDelay(tipd_DI1));
   VitalWireDelay (DI2_ipd, DI2, VitalExtendToFillDelay(tipd_DI2));
   VitalWireDelay (DI3_ipd, DI3, VitalExtendToFillDelay(tipd_DI3));
   VitalWireDelay (DI4_ipd, DI4, VitalExtendToFillDelay(tipd_DI4));
   VitalWireDelay (DI5_ipd, DI5, VitalExtendToFillDelay(tipd_DI5));
   VitalWireDelay (DI6_ipd, DI6, VitalExtendToFillDelay(tipd_DI6));
   VitalWireDelay (DI7_ipd, DI7, VitalExtendToFillDelay(tipd_DI7));
   VitalWireDelay (DI8_ipd, DI8, VitalExtendToFillDelay(tipd_DI8));
   VitalWireDelay (WRB_ipd, WRB, VitalExtendToFillDelay(tipd_WRB));
   VitalWireDelay (RDB_ipd, RDB, VitalExtendToFillDelay(tipd_RDB));
   VitalWireDelay (WBLKB_ipd, WBLKB, VitalExtendToFillDelay(tipd_WBLKB));
   VitalWireDelay (RBLKB_ipd, RBLKB, VitalExtendToFillDelay(tipd_RBLKB));
   VitalWireDelay (PARODD_ipd, PARODD, VitalExtendToFillDelay(tipd_PARODD));
   VitalWireDelay (RESET_ipd, RESET, VitalExtendToFillDelay(tipd_RESET));
   VitalWireDelay (RCLKS_ipd, RCLKS, VitalExtendToFillDelay(tipd_RCLKS));
   VitalWireDelay (WCLKS_ipd, WCLKS, VitalExtendToFillDelay(tipd_WCLKS));
   VitalWireDelay (DIS_ipd, DIS, VitalExtendToFillDelay(tipd_DIS));

   end block WIRE_DELAY;

   ---------------------------------------------------------------
   --                  Behavior Section                         --
   ---------------------------------------------------------------


    WBint       <= ( WRB_ipd or WBLKB_ipd );
    RBint       <= ( RDB_ipd or RBLKB_ipd);

    VITALBehavior : process (
                          LEVEL0_ipd, LEVEL1_ipd, LEVEL2_ipd, LEVEL3_ipd, LEVEL4_ipd, LEVEL5_ipd, LEVEL6_ipd, LEVEL7_ipd, 
                          LGDEP0_ipd, LGDEP1_ipd, LGDEP2_ipd, 
                          DI0_ipd, DI1_ipd, DI2_ipd, DI3_ipd, DI4_ipd, DI5_ipd, DI6_ipd, DI7_ipd, DI8_ipd, 
                          RCLKS_ipd, 
                          WCLKS_ipd, 
                          WBint, RBint, WRB_ipd, WBLKB_ipd, RDB_ipd, RBLKB_ipd , DIS_ipd, PARODD_ipd, RESET_ipd
                          )

     -- some internal veriable declaration
     variable RAM_di_int   : std_logic_vector(8 downto 0);
     variable memory_array : MEM_TYPE  := (others =>(others => 'X'));
     variable do_par       : std_logic := 'X';
     variable tmp_par      : std_logic := 'X';
     variable tmp_par2     : std_logic := 'X';
     variable wpe_var      : std_logic := 'X';
     variable temp         : integer   := 0;
     variable thresh       : integer   := 0;
     variable depth        : integer   := 0;
     variable WADDR        : integer   := 0;
     variable WADDR_wrap   : integer   := 0;
     variable RADDR        : integer   := 0;
     variable RADDR_wrap   : integer   := 0;

     type SL_TO_INT is array(std_ulogic range 'U' to '-') of integer;
     constant INT :SL_TO_INT := (-65, -65, 0, 1, -65, -65, 0, 1, -65);

     --  Read Timing Check Results
     variable PeriodData_RESET           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RESET                : X01                 := '0';
     variable Tviol_PARODD_RCLKS_posedge : X01                 := '0';
     variable TmDt_PARODD_RCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RDB_RCLKS_posedge    : X01                 := '0';
     variable TmDt_RDB_RCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RBLKB_RCLKS_posedge  : X01                 := '0';
     variable TmDt_RBLKB_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_RCLKS_posedge  : X01                 := '0';
     variable Tmkr_RESET_RCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_RCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_RCLKS                : X01                 := '0';
     variable Tviol_DI0_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI0_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI1_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI1_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI2_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI2_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI3_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI3_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI4_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI4_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI5_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI5_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI6_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI6_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI7_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI7_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_DI8_WCLKS_posedge    : X01                 := '0';
     variable TmDt_DI8_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_PARODD_WCLKS_posedge : X01                 := '0';
     variable TmDt_PARODD_WCLKS_posedge  : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WRB_WCLKS_posedge    : X01                 := '0';
     variable TmDt_WRB_WCLKS_posedge     : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_WBLKB_WCLKS_posedge  : X01                 := '0';
     variable TmDt_WBLKB_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable Tviol_RESET_WCLKS_posedge  : X01                 := '0';
     variable Tmkr_RESET_WCLKS_posedge   : VitalTimingDataType := VitalTimingDataInit;
     variable PeriodData_WCLKS           : VitalPeriodDataType := VitalPeriodDataInit;
     variable Pviol_WCLKS                : X01                 := '0';

     -- functional Results


     variable DO0_zd   : std_ulogic;
     variable DO1_zd   : std_ulogic;
     variable DO2_zd   : std_ulogic;
     variable DO3_zd   : std_ulogic;
     variable DO4_zd   : std_ulogic;
     variable DO5_zd   : std_ulogic;
     variable DO6_zd   : std_ulogic;
     variable DO7_zd   : std_ulogic;
     variable DO8_zd   : std_ulogic;
     variable RPE_zd   : std_ulogic;
     variable WPE_zd   : std_ulogic;
     variable DOS_zd   : std_ulogic;
     variable FULL_zd  : std_ulogic;
     variable EMPTY_zd : std_ulogic;
     variable EQTH_zd  : std_ulogic;
     variable GEQTH_zd : std_ulogic;
     variable FULL_tmp  : std_ulogic;
     variable EMPTY_tmp : std_ulogic;
     variable EQTH_tmp  : std_ulogic;
     variable GEQTH_tmp : std_ulogic;

     -- Output Glitch Detection Support Variables
     variable DO0_GlitchData   : VitalGlitchDataType;
     variable DO1_GlitchData   : VitalGlitchDataType;
     variable DO2_GlitchData   : VitalGlitchDataType;
     variable DO3_GlitchData   : VitalGlitchDataType;
     variable DO4_GlitchData   : VitalGlitchDataType;
     variable DO5_GlitchData   : VitalGlitchDataType;
     variable DO6_GlitchData   : VitalGlitchDataType;
     variable DO7_GlitchData   : VitalGlitchDataType;
     variable DO8_GlitchData   : VitalGlitchDataType;
     variable DOS_GlitchData   : VitalGlitchDataType;
     variable FULL_GlitchData  : VitalGlitchDataType;
     variable EMPTY_GlitchData : VitalGlitchDataType;
     variable EQTH_GlitchData  : VitalGlitchDataType;
     variable GEQTH_GlitchData : VitalGlitchDataType;

     -- last value variables
     variable WCLKS_previous   : std_ulogic := 'X';
     variable RCLKS_previous   : std_ulogic := 'X';
     variable RBint_delayed    : std_ulogic := 'X';
     variable RBint_previous   : std_ulogic := 'X';
     variable WBint_delayed    : std_ulogic := 'X';
     variable WBint_previous   : std_ulogic := 'X';
     variable DIS_previous     : std_ulogic := 'X';
     variable RESET_previous   : std_ulogic := 'X';
     variable RESET_delayed    : std_ulogic := 'X';
     variable PARODD_previous  : std_ulogic := 'X';
     variable PARODD_delayed   : std_ulogic := 'X';
     variable DI0_delayed      : std_ulogic := 'X';
     variable DI1_delayed      : std_ulogic := 'X';
     variable DI2_delayed      : std_ulogic := 'X';
     variable DI3_delayed      : std_ulogic := 'X';
     variable DI4_delayed      : std_ulogic := 'X';
     variable DI5_delayed      : std_ulogic := 'X';
     variable DI6_delayed      : std_ulogic := 'X';
     variable DI7_delayed      : std_ulogic := 'X';
     variable DI8_delayed      : std_ulogic := 'X';
     variable DI0_previous     : std_ulogic := 'X';
     variable DI1_previous     : std_ulogic := 'X';
     variable DI2_previous     : std_ulogic := 'X';
     variable DI3_previous     : std_ulogic := 'X';
     variable DI4_previous     : std_ulogic := 'X';
     variable DI5_previous     : std_ulogic := 'X';
     variable DI6_previous     : std_ulogic := 'X';
     variable DI7_previous     : std_ulogic := 'X';
     variable DI8_previous     : std_ulogic := 'X';
     variable LGDEP0_delayed   : std_ulogic := 'X';
     variable LGDEP1_delayed   : std_ulogic := 'X';
     variable LGDEP2_delayed   : std_ulogic := 'X';
     variable LGDEP0_previous  : std_ulogic := 'X';
     variable LGDEP1_previous  : std_ulogic := 'X';
     variable LGDEP2_previous  : std_ulogic := 'X';
     variable LEVEL0_delayed   : std_ulogic := 'X';
     variable LEVEL1_delayed   : std_ulogic := 'X';
     variable LEVEL2_delayed   : std_ulogic := 'X';
     variable LEVEL3_delayed   : std_ulogic := 'X';
     variable LEVEL4_delayed   : std_ulogic := 'X';
     variable LEVEL5_delayed   : std_ulogic := 'X';
     variable LEVEL6_delayed   : std_ulogic := 'X';
     variable LEVEL7_delayed   : std_ulogic := 'X';
     variable LEVEL0_previous  : std_ulogic := 'X';
     variable LEVEL1_previous  : std_ulogic := 'X';
     variable LEVEL2_previous  : std_ulogic := 'X';
     variable LEVEL3_previous  : std_ulogic := 'X';
     variable LEVEL4_previous  : std_ulogic := 'X';
     variable LEVEL5_previous  : std_ulogic := 'X';
     variable LEVEL6_previous  : std_ulogic := 'X';
     variable LEVEL7_previous  : std_ulogic := 'X';

     --  Pipelined temporary results
     variable RPE_stg1         : std_ulogic := 'X';
     variable DO0_stg1         : std_ulogic := 'X';
     variable DO1_stg1         : std_ulogic := 'X';
     variable DO2_stg1         : std_ulogic := 'X';
     variable DO3_stg1         : std_ulogic := 'X';
     variable DO4_stg1         : std_ulogic := 'X';
     variable DO5_stg1         : std_ulogic := 'X';
     variable DO6_stg1         : std_ulogic := 'X';
     variable DO7_stg1         : std_ulogic := 'X';
     variable DO8_stg1         : std_ulogic := 'X';

     -- Special variables to control flags
     variable hold_empty_low   : integer := 0;
     variable hold_eqth_high   : integer := 0;
     variable hold_geqth_high  : integer := 0;
     variable hold_full_low    : integer := 0;
     variable hold_empty_high  : integer := 0;
     variable hold_eqth_low    : integer := 0;
     variable hold_geqth_low   : integer := 0;

     variable WCLKS_re         : Time;
     variable WCLKS_fe         : Time;
     variable WCLKS_fe_prev    : Time;
     variable WB_re            : Time;
     variable RESET_re         : Time;

 begin -- process VITALBehavior

 if (TimingCheckOn) then
   ---------------------------------------------------------
   -- # Read Timing Check Section                         --
   ---------------------------------------------------------

   -- recovery / removal check for RCLKS to RESET signal ;
       VitalRecoveryRemovalCheck ( Tviol_RESET_RCLKS_posedge,
                             Tmkr_RESET_RCLKS_posedge,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             trecovery_RESET_RCLKS_posedge_negedge,
                             thold_RESET_RCLKS_posedge_posedge,
                             TRUE,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'), 
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             TRUE,
                             TRUE,
                             WARNING
                             );

   -- setup hold REN, RBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_RDB_RCLKS_posedge,
                             TmDt_RDB_RCLKS_posedge,
                             RDB_ipd, "RDB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns,
                             tsetup_RDB_RCLKS_posedge_posedge,
                             tsetup_RDB_RCLKS_negedge_posedge,
                             thold_RDB_RCLKS_posedge_posedge,
                             thold_RDB_RCLKS_negedge_posedge,
                             ((TO_X01(RBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_RBLKB_RCLKS_posedge,
                             TmDt_RBLKB_RCLKS_posedge,
                             RBLKB_ipd, "RBLKB",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_RBLKB_RCLKS_posedge_posedge,
                             tsetup_RBLKB_RCLKS_negedge_posedge,
                             thold_RBLKB_RCLKS_posedge_posedge,
                             thold_RBLKB_RCLKS_negedge_posedge,
                             ((TO_X01(RDB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(EMPTY_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_PARODD_RCLKS_posedge,
                             TmDt_PARODD_RCLKS_posedge,
                             PARODD_ipd, "PARODD",
                             0.0 ns,
                             RCLKS_ipd, "RCLKS",
                             0.0 ns, 
                             tsetup_PARODD_RCLKS_posedge_posedge,
                             tsetup_PARODD_RCLKS_negedge_posedge,
                             thold_PARODD_RCLKS_posedge_posedge,
                             thold_PARODD_RCLKS_negedge_posedge,
                             (TO_X01(RESET_ipd) = '1'),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

  --   Period of RCLK
      VitalPeriodPulseCheck ( Pviol_RCLKS,
                              PeriodData_RCLKS,
                              RCLKS_ipd, "RCLKS",
                              0.0 ns,
                              tperiod_RCLKS,
                              tpw_RCLKS_posedge,
                              tpw_RCLKS_negedge,
                              (TO_X01(RDB) = '0') AND (TO_X01(RBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(EMPTY_zd) = '0'),
                              InstancePath & "/FIFO256x9SSRP",
                              True,
                              True,
                              WARNING
                              );
      VitalPeriodPulseCheck ( Pviol_RESET,
                              PeriodData_RESET,
                              RESET_ipd, "RESET",
                              0.0 ns,
                              tpw_RESET_negedge,
                              0.0 ns,
                              tpw_RESET_negedge,
                              True,
                              InstancePath & "/FIFO256x9SSRP",
                              True,
                              True,
                              WARNING
                              );
   ---------------------------------------------------------
   -- # Write Timing Check Section                        --
   ---------------------------------------------------------

       -- recovery / removal check for WCLKS to RESET signal ;
       VitalRecoveryRemovalCheck ( Tviol_RESET_WCLKS_posedge,
                             Tmkr_RESET_WCLKS_posedge,
                             RESET_ipd, "RESET",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns,
                             trecovery_RESET_WCLKS_posedge_negedge,
                             thold_RESET_WCLKS_posedge_posedge,
                             TRUE,
                             (TO_X01(EMPTY_zd) = '1') AND (TO_X01(FULL_zd) = '0'), 
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             TRUE,
                             TRUE,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI0_WCLKS_posedge,
                             TmDt_DI0_WCLKS_posedge,
                             DI0_ipd, "DI0",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI0_WCLKS_posedge_posedge,
                             tsetup_DI0_WCLKS_negedge_posedge,
                             thold_DI0_WCLKS_posedge_posedge,
                             thold_DI0_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI1_WCLKS_posedge,
                             TmDt_DI1_WCLKS_posedge,
                             DI1_ipd, "DI1",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI1_WCLKS_posedge_posedge,
                             tsetup_DI1_WCLKS_negedge_posedge,
                             thold_DI1_WCLKS_posedge_posedge,
                             thold_DI1_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI2_WCLKS_posedge,
                             TmDt_DI2_WCLKS_posedge,
                             DI2_ipd, "DI2",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI2_WCLKS_posedge_posedge,
                             tsetup_DI2_WCLKS_negedge_posedge,
                             thold_DI2_WCLKS_posedge_posedge,
                             thold_DI2_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI3_WCLKS_posedge,
                             TmDt_DI3_WCLKS_posedge,
                             DI3_ipd, "DI3",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI3_WCLKS_posedge_posedge,
                             tsetup_DI3_WCLKS_negedge_posedge,
                             thold_DI3_WCLKS_posedge_posedge,
                             thold_DI3_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI4_WCLKS_posedge,
                             TmDt_DI4_WCLKS_posedge,
                             DI4_ipd, "DI4",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI4_WCLKS_posedge_posedge,
                             tsetup_DI4_WCLKS_negedge_posedge,
                             thold_DI4_WCLKS_posedge_posedge,
                             thold_DI4_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI5_WCLKS_posedge,
                             TmDt_DI5_WCLKS_posedge,
                             DI5_ipd, "DI5",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI5_WCLKS_posedge_posedge,
                             tsetup_DI5_WCLKS_negedge_posedge,
                             thold_DI5_WCLKS_posedge_posedge,
                             thold_DI5_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI6_WCLKS_posedge,
                             TmDt_DI6_WCLKS_posedge,
                             DI6_ipd, "DI6",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI6_WCLKS_posedge_posedge,
                             tsetup_DI6_WCLKS_negedge_posedge,
                             thold_DI6_WCLKS_posedge_posedge,
                             thold_DI6_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI7_WCLKS_posedge,
                             TmDt_DI7_WCLKS_posedge,
                             DI7_ipd, "DI7",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI7_WCLKS_posedge_posedge,
                             tsetup_DI7_WCLKS_negedge_posedge,
                             thold_DI7_WCLKS_posedge_posedge,
                             thold_DI7_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_DI8_WCLKS_posedge,
                             TmDt_DI8_WCLKS_posedge,
                             DI8_ipd, "DI8",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_DI8_WCLKS_posedge_posedge,
                             tsetup_DI8_WCLKS_negedge_posedge,
                             thold_DI8_WCLKS_posedge_posedge,
                             thold_DI8_WCLKS_negedge_posedge,
                             ((TO_X01(WBint) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

   -- setup hold WEN, WBLK low when RCLK rising
       VitalSetupHoldCheck ( Tviol_WRB_WCLKS_posedge,
                             TmDt_WRB_WCLKS_posedge,
                             WRB_ipd, "WRB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WRB_WCLKS_posedge_posedge,
                             tsetup_WRB_WCLKS_negedge_posedge,
                             thold_WRB_WCLKS_posedge_posedge,
                             thold_WRB_WCLKS_negedge_posedge,
                             ((TO_X01(WBLKB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_WBLKB_WCLKS_posedge,
                             TmDt_WBLKB_WCLKS_posedge,
                             WBLKB_ipd, "WBLKB",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_WBLKB_WCLKS_posedge_posedge,
                             tsetup_WBLKB_WCLKS_negedge_posedge,
                             thold_WBLKB_WCLKS_posedge_posedge,
                             thold_WBLKB_WCLKS_negedge_posedge,
                             ((TO_X01(WRB_ipd) = '0') AND (TO_X01(RESET_ipd) = '1') AND (TO_X01(FULL_zd) = '0')),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

       VitalSetupHoldCheck ( Tviol_PARODD_WCLKS_posedge,
                             TmDt_PARODD_WCLKS_posedge,
                             PARODD_ipd, "PARODD",
                             0.0 ns,
                             WCLKS_ipd, "WCLKS",
                             0.0 ns, 
                             tsetup_PARODD_WCLKS_posedge_posedge,
                             tsetup_PARODD_WCLKS_negedge_posedge,
                             thold_PARODD_WCLKS_posedge_posedge,
                             thold_PARODD_WCLKS_negedge_posedge,
                             ((TO_X01(RBint) = '0') AND (TO_X01(RESET_ipd) = '1')),
                             '/',
                             InstancePath & "/FIFO256x9SSRP",
                             True,
                             True,
                             WARNING
                             );

  --   Period of WCLK
      VitalPeriodPulseCheck ( Pviol_WCLKS,
                              PeriodData_WCLKS,
                              WCLKS_ipd, "WCLKS",
                              0.0 ns,
                              tperiod_WCLKS,
                              tpw_WCLKS_posedge,
                              tpw_WCLKS_negedge,
                              (TO_X01(WRB) = '0') AND (TO_X01(WBLKB) = '0') AND (TO_X01(RESET) = '1') AND (TO_X01(FULL_zd) ='0'),
                              InstancePath & "/FIFO256x9SSRP",
                              True,
                              True,
                              WARNING
                              );
 end if;

   ------------------------------------------------------------
   --               FIFO RESET                               --
   ------------------------------------------------------------

   if ( RESET_ipd'event and RESET_ipd = '0' ) then
       WADDR      := 0;
       RADDR      := 0;
       WADDR_wrap := 0;
       RADDR_wrap := 0;
       FULL_tmp   := '0';
       EMPTY_tmp  := '1';
       EQTH_tmp   := '0';
       GEQTH_tmp  := '0';
       WRITE_AT_PREV_EDGE <='0';
       READ_AT_PREV_EDGE <='0';
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
       hold_full_low   := 0;
       hold_empty_high := 0;
       hold_eqth_low   := 0;
       hold_geqth_low  := 0;
   end if;

   if ( WCLKS_ipd'event and WCLKS_ipd = '1' ) then
     WCLKS_re := now;
   end if;
      
   if ( WBint'event and WBint = '1' ) then
     WB_re := now;
   end if;
      
   if ( RESET_ipd'event and RESET_ipd = '1' ) then
     RESET_re := now;
     if ( TO_X01 ( WCLKS_ipd ) = '1' ) then
       if ( WCLKS_re = WB_re ) then
         hold_full_low   := 1; -- until next reset
         hold_empty_high := 1;
         hold_eqth_low   := 1;
         hold_geqth_low  := 1;
       elsif ( TO_X01 ( WBint ) = '0' ) then
         EMPTY_zd        := '0';
         EQTH_zd         := '1';
         GEQTH_zd        := '1';
         hold_empty_low  := 1; -- until next WCLKS falling edge
         hold_eqth_high  := 1;
         hold_geqth_high := 1;
       elsif ( WCLKS_re < WB_re ) then
         EMPTY_zd        := '0';
         EQTH_zd         := '1';
         GEQTH_zd        := '1';
         hold_empty_low  := 1; -- until next WCLKS falling edge
         hold_eqth_high  := 1;
         hold_geqth_high := 1;
       elsif ( WB_re < WCLKS_re ) then
         hold_empty_low  := 0; -- expected behavior
         hold_eqth_high  := 0;
         hold_geqth_high := 0;
         hold_full_low   := 0;
         hold_empty_high := 0;
         hold_eqth_low   := 0;
         hold_geqth_low  := 0;
       end if;
     else
       hold_empty_low  := 0; -- expected behavior
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
       hold_full_low   := 0;
       hold_empty_high := 0;
       hold_eqth_low   := 0;
       hold_geqth_low  := 0;
     end if;
   end if;

   if ( WCLKS_ipd'event and WCLKS_ipd = '0' ) then
     WCLKS_fe_prev := WCLKS_fe;
     WCLKS_fe := now;
     if (( TO_X01 ( RESET_ipd ) = '1' ) and ( WCLKS_fe_prev < RESET_re )) then
       hold_empty_low  := 0;
       hold_eqth_high  := 0;
       hold_geqth_high := 0;
     end if;
   end if;


   ------------------------------------------------------------
   --         WPE generating block                            -
   ------------------------------------------------------------

    if (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') then
      tmp_par  := DI7_ipd XOR DI6_ipd XOR DI5_ipd XOR DI4_ipd XOR DI3_ipd XOR DI2_ipd XOR DI1_ipd XOR DI0_ipd;
      par_f  <= tmp_par ;
      if (tmp_par /= PARODD_ipd) then
        wpe_var  :=  '1';
      else
        wpe_var  :=  '0';
      end if;
      RAM_di_int(8) := wpe_var;
      WPE_zd := wpe_var;
    end if;

   -----------------------------------------------------------
   --     DOS signal                                        --
   -----------------------------------------------------------

   if(DIS_ipd'event)  then
      DOS_zd := DIS_ipd;
   end if; 

   -----------------------------------------------------------
   --    calculate the depth and levels                     --
   -----------------------------------------------------------

    temp :=((INT(LGDEP2_delayed)*4) + (INT(LGDEP1_delayed)*2) + 
           (INT(LGDEP0_delayed)*1));

    case temp is 
         when 0 => depth := 2;
         when 1 => depth := 4;
         when 2 => depth := 8;
         when 3 => depth := 16;
         when 4 => depth := 32;
         when 5 => depth := 64;
         when 6 => depth := 128;
         when 7 => depth := 256;
         when others => depth := 0;
    end case;

    -- thresh value

    thresh := (INT(LEVEL7_delayed)*128) + (INT(LEVEL6_delayed)*64) + 
               (INT(LEVEL5_delayed)*32) + (INT(LEVEL4_delayed)*16) + 
               (INT(LEVEL3_delayed)*8) + (INT(LEVEL2_delayed)*4) + 
               (INT(LEVEL1_delayed)*2) + (INT(LEVEL0_delayed)*1); 

    if ( thresh = 0 or thresh = 255 ) then
      assert false
        report " Illegal level configuration, LEVEL cannot be 0 or 255 "
        severity failure;
    end if;

   ------------------------------------------------------------
   -- # Write Functional Section                             --
   ------------------------------------------------------------

   if(TO_X01(WCLKS_ipd)='X') then
    if(RESET_delayed = '1') then
     if (WBint_delayed = '0') then
      if (TO_X01(WCLKS_previous) /= 'X') then
        assert false
        report ": WCLK unknown"
        severity Error;
      end if;
     end if;
    end if;
   elsif (WCLKS_ipd'EVENT AND WCLKS_ipd = '1') AND (TO_X01(RESET_ipd) = '1')then
     WRITE_AT_PREV_EDGE <='0';
     case (TO_X01(WBint_delayed)) is 
      when '1' =>
                null;
      when '0' => 
         if(FULL_zd = '0') then 
         RAM_di_int(7 downto 0) := DI7_delayed & DI6_delayed & DI5_delayed & 
                                    DI4_delayed & DI3_delayed & DI2_delayed & 
                                    DI1_delayed & DI0_delayed;
         memory_array(WADDR) := RAM_di_int;
         WRITE_AT_PREV_EDGE <='1';
         if(WADDR <depth-1  ) then
           WADDR := WADDR + 1;
         elsif( WADDR  = depth-1) then
           WADDR := 0;
           WADDR_wrap := 1 - WADDR_wrap;
         end if;
        end if;
       when others => 
        if (TO_X01(WBint_previous) /= 'X') then
          assert false
          report ": WBLKB or WRB unknown"
          severity Error;
          end if;
        end case;
     elsif(WCLKS_ipd'EVENT AND WCLKS_ipd = '0')  AND (TO_X01(RESET_delayed) = '1') AND (TO_X01(WRITE_AT_PREV_EDGE) = '1')then
        WRITE_AT_PREV_EDGE <='0';
        if(WADDR   = RADDR ) then
         if(RADDR_wrap /= WADDR_wrap) then
          FULL_tmp := '1';
          EMPTY_tmp :='0';
         end if;
        end if;
        if(WADDR   /= RADDR ) then
          EMPTY_tmp := '0';
        end if;
          if(RADDR_wrap = WADDR_wrap) then
            if(WADDR - RADDR = thresh ) then
               EQTH_tmp := '1';
            else 
               EQTH_tmp := '0';
            end if;
            if(WADDR - RADDR >= thresh ) then
                GEQTH_tmp := '1';
            else 
                GEQTH_tmp := '0';
            end if;
          else 
           if((depth -RADDR + WADDR) = thresh ) then
               EQTH_tmp := '1';
            else 
               EQTH_tmp := '0';
            end if;
            if((depth -RADDR + WADDR) >= thresh ) then
                GEQTH_tmp := '1';
            else 
                GEQTH_tmp := '0';
            end if;
           end if; 
      else
       null;
    end if;


  --------------------------------------------------------------------
  --          FIFO READ SECTION........                             --
  --------------------------------------------------------------------

  if (TO_X01(RCLKS_ipd)='X') then
    if(RESET_ipd /= '0') then
    if(TO_X01(RBint_delayed) /= '1') then
      if(TO_X01(RCLKS_previous) /= 'X') then
        assert false
        report ": RCLK unknown"
        severity Error;
        DO0_zd  := 'X';
        DO1_zd  := 'X';
        DO2_zd  := 'X';
        DO3_zd  := 'X';
        DO4_zd  := 'X';
        DO5_zd  := 'X';
        DO6_zd  := 'X';
        DO7_zd  := 'X';
        DO8_zd  := 'X';
      end if;
     end if;
    end if;
   elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='1') AND (TO_X01(RESET_delayed) = '1')) then
     DO0_zd := DO0_stg1;
     DO1_zd := DO1_stg1;
     DO2_zd := DO2_stg1;
     DO3_zd := DO3_stg1;
     DO4_zd := DO4_stg1;
     DO5_zd := DO5_stg1;
     DO6_zd := DO6_stg1;
     DO7_zd := DO7_stg1;
     DO8_zd := DO8_stg1;
     RPE_zd := RPE_stg1;
     READ_AT_PREV_EDGE <='0';
     case (TO_X01(RBint_delayed)) is
        when '1' =>
                null;
        when '0' =>
         if(TO_X01(EMPTY_zd) /= '1') then 
           DO0_stg1  := memory_array(RADDR)(0);
           DO1_stg1  := memory_array(RADDR)(1);
           DO2_stg1  := memory_array(RADDR)(2);
           DO3_stg1  := memory_array(RADDR)(3);
           DO4_stg1  := memory_array(RADDR)(4);
           DO5_stg1  := memory_array(RADDR)(5);
           DO6_stg1  := memory_array(RADDR)(6);
           DO7_stg1  := memory_array(RADDR)(7);
           DO8_stg1  := memory_array(RADDR)(8);
           READ_AT_PREV_EDGE <='1';
           if(RADDR <depth-1  ) then
             RADDR := RADDR + 1;
           else
             RADDR :=(RADDR +1) mod  depth;
             RADDR_wrap :=1 - RADDR_wrap;
           end if;
      do_par  := DO8_stg1 XOR DO7_stg1 XOR DO6_stg1 XOR DO5_stg1 XOR DO4_stg1 XOR DO3_stg1 XOR
                 DO2_stg1 XOR DO1_stg1 XOR DO0_stg1;
            par_f <= do_par;
            if (do_par = 'X') then
             RPE_stg1 := 'X';
            elsif (do_par /= PARODD_delayed) then
             RPE_stg1  :=  '1';
            else
             RPE_stg1  :=  '0';
            end if;
         end if;
     when others =>
       if (TO_X01(RBint_previous) /= 'X') then
        assert false
        report ": RDB or RBLKB unknown"
        severity Error;
        end if;
           DO0_stg1  := 'X';
           DO1_stg1  := 'X';
           DO2_stg1  := 'X';
           DO3_stg1  := 'X';
           DO4_stg1  := 'X';
           DO5_stg1  := 'X';
           DO6_stg1  := 'X';
           DO7_stg1  := 'X';
           DO8_stg1  := 'X';
     end case;
  elsif (RCLKS_ipd'event and (TO_X01(RCLKS_ipd)='0') AND (TO_X01(RESET_delayed) = '1') AND (TO_X01(READ_AT_PREV_EDGE) = '1')) then
   READ_AT_PREV_EDGE <='0';
   if(RADDR = WADDR ) then
    if(RADDR_wrap = WADDR_wrap) then
       EMPTY_tmp := '1';
       FULL_tmp  := '0';
    end if;
   end if;
   if(RADDR /= WADDR ) then
    FULL_tmp  := '0';
   end if;
    if(WADDR_wrap = RADDR_wrap ) then
     if((WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((WADDR - RADDR) >= thresh  ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    else 
     if((depth + WADDR - RADDR) = thresh ) then
       EQTH_tmp := '1';
     else
       EQTH_tmp := '0';
     end if;
     if((depth + WADDR - RADDR) >= thresh ) then
       GEQTH_tmp := '1';
     else
       GEQTH_tmp := '0';
     end if;
    end if;
 else 
    null;
 end if;

   -- Mimic odd silicon flag behavior coming out of RESET with WB low
   
   if ( hold_full_low = 1 ) then
     FULL_zd := '0';
   else
     FULL_zd := FULL_tmp;
   end if;

   if ( hold_empty_low = 1 ) then
     EMPTY_zd := '0';
   elsif ( hold_empty_high = 1 ) then
     EMPTY_zd := '1';
   else
     EMPTY_zd := EMPTY_tmp;
   end if;

   if ( hold_eqth_high = 1 ) then
     EQTH_zd := '1';
   elsif ( hold_eqth_low = 1 ) then
     EQTH_zd := '0';
   else
     EQTH_zd := EQTH_tmp;
   end if;

   -- If LEVEL greater than DEPTH then GEQTH mimics FULL
   
   if ( hold_geqth_high = 1 ) then
     GEQTH_zd := '1';
   elsif ( hold_geqth_low = 1 ) then
     GEQTH_zd := '0';
   else
     if ( thresh > depth ) then
       GEQTH_zd := FULL_zd;
     else
       GEQTH_zd := GEQTH_tmp;
     end if;
   end if;


  -------------------------------------------------------------------
  --         Internal variable assignment section                  --
  -------------------------------------------------------------------

       WCLKS_previous  := WCLKS_ipd;
       RCLKS_previous   := RCLKS_ipd;
       RBint_previous   := RBint_delayed;
       RBint_delayed    := RBint;
       WBint_previous   := WBint_delayed;
       WBint_delayed    := WBint;
       DI0_delayed      := DI0_ipd;
       DI1_delayed      := DI1_ipd;
       DI2_delayed      := DI2_ipd;
       DI3_delayed      := DI3_ipd;
       DI4_delayed      := DI4_ipd;
       DI5_delayed      := DI5_ipd;
       DI6_delayed      := DI6_ipd;
       DI7_delayed      := DI7_ipd;
       DI8_delayed      := DI8_ipd;
       LGDEP0_previous  := LGDEP0_delayed;
       LGDEP0_delayed   := LGDEP0_ipd;
       LGDEP1_previous  := LGDEP1_delayed;
       LGDEP1_delayed   := LGDEP1_ipd;
       LGDEP2_previous  := LGDEP2_delayed;
       LGDEP2_delayed   := LGDEP2_ipd;
       LEVEL0_previous  := LEVEL0_delayed;
       LEVEL0_delayed   := LEVEL0_ipd;
       LEVEL1_previous  := LEVEL1_delayed;
       LEVEL1_delayed   := LEVEL1_ipd;
       LEVEL2_previous  := LEVEL2_delayed;
       LEVEL2_delayed   := LEVEL2_ipd;
       LEVEL3_previous  := LEVEL3_delayed;
       LEVEL3_delayed   := LEVEL3_ipd;
       LEVEL4_previous  := LEVEL4_delayed;
       LEVEL4_delayed   := LEVEL4_ipd;
       LEVEL5_previous  := LEVEL5_delayed;
       LEVEL5_delayed   := LEVEL5_ipd;
       LEVEL6_previous  := LEVEL6_delayed;
       LEVEL6_delayed   := LEVEL6_ipd;
       LEVEL7_previous  := LEVEL7_delayed;
       LEVEL7_delayed   := LEVEL7_ipd;
       PARODD_previous  := PARODD_delayed; 
       PARODD_delayed   := PARODD_ipd;
       RESET_previous   := RESET_delayed; 
       RESET_delayed    := RESET_ipd;


 -------------------------------------------------------------
 --              Path Delay Section                         --
 -------------------------------------------------------------

     VitalPathDelay01Z (
             OutSignal     => DOS,
             GlitchData    => DOS_GlitchData,
             OutSignalName => "DOS",
             OutTemp       => DOS_zd,

             Paths =>   (0 => (DIS_ipd'last_event,
                                VitalExtendToFillDelay(tpd_DIS_DOS), true)),

             DefaultDelay  => VitalZeroDelay01Z,
             Mode          => Onevent,
             Xon           => Xon,
             MsgOn         => MsgOn,
             MsgSeverity   => WARNING
             );

     VitalPathDelay01Z (
           OutSignal     => DO0,
           GlitchData    => DO0_GlitchData,
           OutSignalName => "DO0",
           OutTemp       => DO0_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO0), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO0), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO1,
           GlitchData    => DO1_GlitchData,
           OutSignalName => "DO1",
           OutTemp       => DO1_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO1), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO1), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO2,
           GlitchData    => DO2_GlitchData,
           OutSignalName => "DO2",
           OutTemp       => DO2_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO2), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO2), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO3,
           GlitchData    => DO3_GlitchData,
           OutSignalName => "DO3",
           OutTemp       => DO3_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO3), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO3), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO4,
           GlitchData    => DO4_GlitchData,
           OutSignalName => "DO4",
           OutTemp       => DO4_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO4), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO4), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO5,
           GlitchData    => DO5_GlitchData,
           OutSignalName => "DO5",
           OutTemp       => DO5_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO5), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO5), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO6,
           GlitchData    => DO6_GlitchData,
           OutSignalName => "DO6",
           OutTemp       => DO6_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO6), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO6), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO7,
           GlitchData    => DO7_GlitchData,
           OutSignalName => "DO7",
           OutTemp       => DO7_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO7), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO7), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => DO8,
           GlitchData    => DO8_GlitchData,
           OutSignalName => "DO8",
           OutTemp       => DO8_zd,

           Paths =>   (0 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_DO8), true),
                       1 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_DO8), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
        );

     VitalPathDelay01Z (
           OutSignal     => FULL,
           GlitchData    => FULL_GlitchData,
           OutSignalName => "FULL",
           OutTemp       => FULL_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_FULL), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_FULL), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_FULL), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EMPTY,
           GlitchData    => EMPTY_GlitchData,
           OutSignalName => "EMPTY",
           OutTemp       => EMPTY_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EMPTY), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_EMPTY), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EMPTY), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => True,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => EQTH,
           GlitchData    => EQTH_GlitchData,
           OutSignalName => "EQTH",
           OutTemp       => EQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_EQTH), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_EQTH), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_EQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );

     VitalPathDelay01Z (
           OutSignal     => GEQTH,
           GlitchData    => GEQTH_GlitchData,
           OutSignalName => "GEQTH",
           OutTemp       => GEQTH_zd,

           Paths =>   (0 => (RESET_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RESET_GEQTH), true),
                       1 => (WCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_WCLKS_GEQTH), true),
                       2 => (RCLKS_ipd'last_event,
                               VitalExtendToFillDelay(tpd_RCLKS_GEQTH), true)),

           DefaultDelay  => VitalZeroDelay01Z,
           Mode          => Onevent,
           Xon           => Xon,
           MsgOn         => MsgOn,
           MsgSeverity   => WARNING
           );


   end process VITALBehavior;

  end VITAL_ACT;
