* BEGIN MODEL LMH6550
*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Corporation.
* Models developed and under copyright by:
* National Semiconductor, Corporation.
*/////////////////////////////////////////////////////////////////////
* Legal Notice:
* The model may be copied, and distributed without any modifications;
* however, reselling or licensing the material is illegal.
* We reserve the right to make changes to the model without prior notice.
* Pspice Models are provided "AS IS, WITH NO WARRANTY OF ANY KIND"
*////////////////////////////////////////////////////////////////////
*////////////////////////////////////////////////////////////////////
* For more information, and our latest models,
* please visit the models section of our website at
*       http://www.national.com/models/
*////////////////////////////////////////////////////////////////////
*MODEL FEATURES INCLUDE OUTPUT SWING, OUTPUT CURRENT
*THRU THE SUPPLIES, GAIN AND PHASE, CLOSED LOOP BANDWIDTH,
*SLEW RATE, COMMON MODE REJECTION WITH FREQUENCY EFFECTS,
*POWER SUPPLY REJECTION, INPUT VOLTAGE NOISE WITH 1/F,
*INPUT CURRENT NOISE, INPUT BIAS CURRENT WITH TEMPCO,
*INPUT OFFSET AND TEMPCO, VCM INPUT OFFSET AND TEMPCO,
*ENABLE WITH ON AND OFF DELAYS, OUTPUT IMPEDANCE, CLOAD
*EFFECTS, VCM SLEW RATE, BALLANCE ERROR VS FREQUENCY,
*OUTPUT SHORT CIRCUIT CURRENT, AND QUIESCENT SUPPLY CURRENT.
*///MODEL TEMP RANGE IS -40 TO +85 DEG C.///
*//////////////////////////////////////////////////////////
* PINOUT ORDER +IN -IN V+ V- +OUT -OUT VCM EN
* PINOUT ORDER  8   1  3  6   4    5    2  7
.SUBCKT LMH6550 8 1 3 6 4 5 2 7
*
Q62 183 183 185 QP
Q63 186 182 183 QP
R70 185 3 2E3
Q64 186 103 187 Q
R71 6 187 2E3
Q65 103 103 188 Q
Q66 3 186 103 Q
R72 6 188 2E3
Q67 189 103 190 Q
R73 6 190 1960
Q68 104 104 191 QP
Q5 6 117 116 QP
R7 118 117 40
Q6 6 119 115 QP 2
Q7 3 112 118 Q 2
Q8 118 102 120 Q 2
R8 6 120 250
Q9 119 102 121 Q 2
R9 6 121 250
Q17 124 104 130 QP 4
Q18 127 103 131 Q 4
R16 6 131 492
C1 115 101 0.83E-12
C2 118 102 0.83E-12
Q19 3 132 133 Q
Q20 134 105 135 QP 2
R17 135 3 252
Q21 136 105 137 QP 2
R18 137 3 250
Q22 105 105 138 QP
R19 138 3 500
R20 134 132 40
R21 5 133 2
R22 139 5 2
Q23 6 140 139 QP
R23 141 140 40
Q24 6 142 134 QP 2
Q25 3 136 141 Q 2
Q26 141 106 143 Q 2
R24 6 143 250
Q27 142 106 144 Q 2
R25 6 144 250
Q28 106 106 145 Q
R26 6 145 500
R27 142 136 24
Q35 147 104 155 QP 4
Q36 150 103 156 Q 4
R32 6 156 492
C3 134 105 0.83E-12
C4 141 106 0.83E-12
R33 149 126 200
R34 110 3 585
Q37 105 157 158 Q
Q38 159 159 160 QP
R36 160 3 800
R37 2 3 60E3
Q39 106 157 109 QP
Q40 161 162 109 QP 2
R58 169 7 6E3
R59 7 3 20E3
Q1 3 107 108 Q
Q2 109 104 110 QP 2
R1 111 3 252
Q3 112 101 113 QP 2
R2 113 3 250
Q4 101 101 114 QP
R3 114 3 500
R4 115 107 40
R5 4 108 2
R6 116 4 2
R69 6 180 5.4E3
Q51 6 169 172 QP
Q52 172 173 174 QP
R60 174 3 1E3
R61 175 3 1E3
Q53 173 173 175 QP
R62 176 173 15.8E3
R63 168 3 33.5E3
Q54 176 177 178 Q
R64 6 171 8E3
R65 6 178 250
Q55 170 170 177 Q 2
Q56 179 170 180 Q
Q57 177 180 6 Q
Q29 6 146 147 QP
Q30 105 148 149 Q
R28 148 147 40
Q31 3 146 150 Q
R38 163 162 200
R39 163 4 2.5003E3
R40 5 163 2.5E3
R41 2 157 200
Q41 102 164 109 QP
Q42 101 164 158 Q
R42 164 2 200
Q43 159 165 158 Q 2
Q44 161 161 166 Q
R43 6 166 800
Q45 158 103 167 Q 2
R44 6 167 500
R45 6 2 60E3
R46 165 163 200
Q46 115 101 111 QP 2
Q49 6 168 169 QP
Q50 168 170 171 Q
Q32 106 151 149 QP
R29 151 150 40
Q33 6 152 153 QP 1.01
R30 154 3 492
R31 155 3 492
Q34 153 104 154 QP 4
Q58 180 177 181 Q 2
R66 170 3 84E3
Q59 3 176 179 Q
Q60 182 172 179 Q
Q61 182 183 184 QP
R67 184 3 2E3
R68 6 181 1150
R74 191 3 2E3
Q69 189 104 192 QP
R75 192 3 2E3
Q70 6 189 104 QP
C5 170 6 0.5E-12
I1 146 152 1.2E-6
I2 123 8 1.2E-6
E2 146 0 153 0 0.99986
V33 152 1 -100E-6
Q10 102 102 122 Q
R10 6 122 500
R11 119 112 24
Q11 6 123 124 QP
Q12 101 125 126 Q
R12 125 124 40
Q13 3 123 127 Q
Q14 102 128 126 QP
R13 128 127 40
Q15 6 8 123 QP
R14 129 3 492
R15 130 3 492
Q16 123 104 129 QP 4
.MODEL Q NPN BF=179.3 VAF=68 RB=80 KF=1E-16 IKF=0.1
.MODEL QP PNP BF=105.95 VAF=68 RB=80 KF=1E-16 IKF=0.1
.ENDS
* END MODEL LMH6550

