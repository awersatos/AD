* BEGIN MODEL LMP8270
* Rev B 5/22/06
*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Corporation.
* Models developed and under copyright by:
* National Semiconductor, Corporation.
*/////////////////////////////////////////////////////////////////////
* Legal Notice:
* The model may be copied, and distributed without any modifications;
* however, reselling or licensing the material is illegal.
* We reserve the right to make changes to the model without prior notice.
* Pspice Models are provided "AS IS, WITH NO WARRANTY OF ANY KIND"
*////////////////////////////////////////////////////////////////////
* For more information, and our latest models,
* please visit the models section of our website at
*       http://www.national.com/models/
*////////////////////////////////////////////////////////////////////
*
* PINOUT ORDER -IN GND A1 A2 OUT VS +IN
* PINOUT ORDER  1   2   3  4  5   6   8
.SUBCKT LMP8270 1 2 3 4 5 6 8
Q20 9 10 11 QON
R10 10 12 100
R11 13 14 100
R12 14 6 20
R13 2 12 20
R16 15 16 2E3
R17 17 18 20
R18 11 19 20
D5 20 6 DD
D6 2 20 DD
D7 21 11 DIN
D8 22 11 DIN
I8 11 21 0.1E-3
I9 11 22 0.1E-3
E3 18 0 6 0 1
D9 23 11 DVN
D10 24 11 DVN
I10 11 23 0.4E-6
I11 11 24 0.4E-6
E4 25 26 23 24 63
G2 27 26 21 22 2.9E-7
E5 28 11 18 11 1
E6 29 11 11 11 1
R30 28 30 1E6
R31 29 31 1E6
R33 11 30 100
R34 11 31 100
C6 28 30 0.2E-12
C7 29 31 0.2E-12
E11 32 33 31 11 0.031
E12 27 32 30 11 0.13
E14 34 11 18 11 0.5
D11 15 18 DD
D12 11 15 DD
M1 35 36 12 12 NOUT L=3U W=200U
M2 37 38 14 14 POUT L=3U W=200U
M3 39 39 17 17 POUT L=3U W=200U
M4 40 41 42 42 PIN L=3U W=22U
M5 43 25 42 42 PIN L=3U W=22U
M8 44 44 19 19 NOUT L=3U W=200U
R43 45 38 100
R44 46 36 100
G3 15 34 47 34 0.2E-3
R45 34 15 6E6
C12 16 20 33E-12
R46 11 40 2.05E3
R47 11 43 2.05E3
C13 40 43 30E-12
C14 27 11 1.5E-12
C15 25 11 1.5E-12
C16 20 0 1E-12
D13 36 9 DD
D14 48 38 DD
Q15 48 13 18 QOP
V18 27 41 -0.35E-3
M16 49 50 51 51 NIN L=3U W=22U
M17 52 25 51 51 NIN L=3U W=22U
R55 49 18 2.05E3
R56 52 18 2.05E3
C20 49 52 30E-12
V19 41 50 0
M18 53 54 55 55 PIN L=6U W=500U
M19 56 57 18 18 PIN L=6U W=500U
V20 18 54 1.9
M21 51 53 11 11 NIN L=6U W=500U
M22 53 53 11 11 NIN L=6U W=500U
G6 15 34 58 34 0.2E-3
I14 39 44 80E-6
M23 57 57 18 18 PIN L=6U W=500U
I15 57 11 100E-6
V21 56 42 0
R59 20 37 50
R60 35 59 50
J1 18 27 18 JC
J2 18 25 18 JC
J3 25 11 25 JC
J4 27 11 27 JC
C21 27 25 0.5E-12
E19 60 34 52 49 1
R61 60 58 10E3
C22 58 34 11E-12
E20 61 34 43 40 1
R62 61 47 10E3
C23 47 34 11E-12
G7 62 34 15 34 -1E-3
G8 34 63 15 34 1E-3
G9 34 64 44 11 1E-3
G10 65 34 18 39 1E-3
D17 65 62 DD
D18 63 64 DD
R66 62 65 100E6
R67 64 63 100E6
R68 65 18 1E3
R69 11 64 1E3
E23 18 45 18 65 1
E24 46 11 64 11 1
R70 63 34 1E6
R71 64 34 1E6
R72 34 65 1E6
R73 34 62 1E6
R77 33 32 1E9
R78 32 27 1E9
R79 26 25 1E9
R80 45 18 1E9
R81 11 46 1E9
R82 34 47 1E9
R83 34 58 1E9
R85 55 56 6.5E3
R86 2 6 1E6
G12 6 2 66 2 -290E-12
I22 2 67 1E-3
D20 67 2 DD
V24 67 66 0.71
R87 2 66 1E6
I23 6 2 618E-6
Q21 68 69 70 QON
R88 69 71 100
R89 72 73 100
R90 73 6 20
R91 2 71 20
R92 74 75 5E3
R93 76 77 20
R94 70 78 20
D22 2 5 DD
D23 79 70 DIN
D24 80 70 DIN
I24 70 79 0.1E-3
I25 70 80 0.1E-3
E26 77 0 6 0 1
D25 81 70 DVN
D26 82 70 DVN
I26 70 81 0.4E-6
I27 70 82 0.4E-6
E27 83 84 81 82 13
G13 4 84 79 80 2.9E-7
E34 85 70 77 70 0.5
D27 74 77 DD
D28 70 74 DD
M24 86 87 71 71 NOUT L=3U W=200U
M25 88 89 73 73 POUT L=3U W=200U
M26 90 90 76 76 POUT L=3U W=200U
M27 91 92 93 93 PIN L=3U W=60U
M28 94 83 93 93 PIN L=3U W=60U
M29 95 95 78 78 NOUT L=3U W=200U
R103 96 89 100
R104 97 87 100
G14 74 85 98 85 0.2E-3
R105 85 74 6E6
C27 75 5 24E-12
R106 70 91 2.05E3
R107 70 94 2.05E3
C28 91 94 30E-12
C29 4 70 4.5E-12
C30 83 70 4.5E-12
C31 5 0 1E-12
D29 87 68 DD
D30 99 89 DD
Q22 99 72 77 QOP
V25 4 92 0
M30 100 101 102 102 NIN L=3U W=60U
M31 103 83 102 102 NIN L=3U W=60U
R108 100 77 2.05E3
R109 103 77 2.05E3
C32 100 103 30E-12
V26 92 101 0
M32 104 105 106 106 PIN L=6U W=500U
M33 107 108 77 77 PIN L=6U W=500U
V27 77 105 1.9
M34 102 104 70 70 NIN L=6U W=500U
M35 104 104 70 70 NIN L=6U W=500U
G15 74 85 109 85 0.2E-3
I28 90 95 80E-6
M36 108 108 77 77 PIN L=6U W=500U
I29 108 70 45E-6
V28 107 93 0
R110 5 88 25
R111 86 110 25
J5 77 4 77 JC
J6 77 83 77 JC
J7 83 70 83 JC
J8 4 70 4 JC
C33 4 83 3.5E-12
E37 111 85 103 100 1
R112 111 109 10E3
C34 109 85 11E-12
E38 112 85 94 91 1
R113 112 98 10E3
C35 98 85 11E-12
G16 113 85 74 85 -1E-3
G17 85 114 74 85 1E-3
G18 85 115 95 70 1E-3
G19 116 85 77 90 1E-3
D31 116 113 DD
D32 114 115 DD
R114 113 116 100E6
R115 115 114 100E6
R116 116 77 1E3
R117 70 115 1E3
E39 77 96 77 116 1
E40 97 70 115 70 1
R118 114 85 1E6
R119 115 85 1E6
R120 85 116 1E6
R121 85 113 1E6
R125 84 83 1E9
R126 96 77 1E9
R127 70 97 1E9
R128 85 98 1E9
R129 85 109 1E9
R131 106 107 6.5E3
D33 5 6 DD
E41 117 70 8 70 1
R132 118 8 200E3
R133 1 118 200E3
E42 119 70 1 70 1
R134 120 117 1E3
R135 119 120 1E3
E44 121 122 8 1 10
V31 122 123 0.5
E45 123 70 124 70 1
R136 124 118 10E3
C72 118 124 1E-9
M37 125 118 70 70 MCP L=3U W=300U
M38 125 126 70 70 MCN L=3U W=300U
E46 126 70 118 70 -1
R137 125 127 1
R138 128 124 10
M39 129 118 70 70 MCMRP L=3U W=300U
M40 129 130 70 70 MCMRN L=3U W=300U
E47 130 70 118 70 -1
V32 131 70 5
R139 129 131 10E3
M41 128 129 70 70 MCMRS L=3U W=3000U
R140 70 124 100
R141 26 20 100E3
R142 132 26 100E3
R143 20 3 100E3
C73 3 0 0.1E-12
R144 70 84 100E3
R145 84 133 50E3
V33 134 122 -0.5
R147 121 127 9E3
C74 26 20 11.4E-12
E48 133 0 5 0 1
E49 118 70 120 70 1
C75 8 118 1E-12
C76 118 1 1E-12
C77 8 70 1E-12
C78 1 70 1E-12
G21 8 70 118 70 4.9E-6
G22 1 70 118 70 4.9E-6
I31 70 135 1E-3
D35 135 70 DD
V37 135 136 0.71
R149 70 136 1E6
E50 132 122 136 70 0.085
E51 137 127 147 134 0.025E-6
R153 147 84 100E3
R154 33 137 92E3
R155 11 33 200E3
R156 147 33 200E3
C79 84 133 25E-12
R157 0 134 1E11
I32 20 2 100E-6
I33 5 2 100E-6
V39 20 59 5E-3
V40 5 110 5E-3
E52 70 0 2 0 1
E53 11 0 2 0 1
RSIN 147 0 1
.MODEL MCP NMOS KP=200U VTO=36.5
.MODEL MCN NMOS KP=200U VTO=2.2
.MODEL MCMRP NMOS KP=200U VTO=27.2
.MODEL MCMRN NMOS KP=200U VTO=2
.MODEL MCMRS NMOS KP=200U VTO=1
.MODEL DD D
.MODEL QON NPN
.MODEL QOP PNP
.MODEL JC NJF
.MODEL DVN D KF=1E-17 IS=1E-16
.MODEL DIN D
.MODEL POUT PMOS KP=200U VTO=-0.7 LAMBDA=0.01
.MODEL NOUT NMOS KP=200U VTO=0.7 LAMBDA=0.01
.MODEL PIN PMOS KP=200U VTO=-0.7
.MODEL NIN NMOS KP=200U VTO=0.7
.MODEL PSW PMOS KP=200U VTO=-0.5 IS=1E-18
.MODEL NSW NMOS KP=200U VTO=0.5 IS=1E-18
.ENDS
* END MODEL LMP8270

