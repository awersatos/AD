*Default PNP Darlington Transistor pkg:TO-92B 1,2,3
*PNP Trans Pinout: C,B,E
.SUBCKT PNP1 1 2 3
Q1 1 2 4 QMOD .1
Q2 1 4 3 QMOD
.MODEL QMOD PNP ()
.ENDS PNP1