--
--                          "num_std.vhd"
--
-- This file contains no vhdl code, this file allows a GUI to reference
-- the pre-compiled file "num_std.mm0" as num_std.vhd.
-- 
-- "num_std.mm0" contains an implementation of the package NUMERIC_STD, this
-- package is part if IEEE Standard 1076.3 "Standard VHDL Synthesis Packages".
--
-- The file "num_bit.mm0" contains the 1076.3 NUMERIC_BIT package.
--
-- Source code for 1076.3 is copyright IEEE and is available from the IEEE.
--
