*//////////////////////////////////////////////////////////////////////
* (C) National Semiconductor, Corporation.
* Models developed and under copyright by:
* National Semiconductor, Corporation.
*/////////////////////////////////////////////////////////////////////
* Legal Notice:
* The model may be copied, and distributed without any modifications;
* however, reselling or licensing the material is illegal.
* We reserve the right to make changes to the model without prior notice.
* Pspice Models are provided "AS IS, WITH NO WARRANTY OF ANY KIND"
*////////////////////////////////////////////////////////////////////
* For more information, and our latest models,
* please visit the models section of our website at
*       http://www.national.com/models/
*////////////////////////////////////////////////////////////////////
* The model below is the CLC5523 renamed as LMH6505 (The LMH6505 is a replacement for the CLC5523 and LMH6504)
* This model simulates the behavior of the LMH6505 for +/-5V supplies only
* LMH6505 SPICE MODEL
* PINOUT ORDER VG VIN RG GND V- OUT I- V+
*
.SUBCKT LMH6505 1 2 63 64 65 66 7 68
*
LP3 3 63 1.0E-9
RLP3 3 63 7.0
LP4 4 64 1.2E-9
RLP4 4 64 7.0
LP5 5 65 1.2E-9
RLP5 5 65 7.0
LP6 6 66 1.0E-9
RLP6 6 66 7.0
LP8 8 68 1.2E-9
RLP8 8 68 7.0
CP27 2 7 0.25E-12
CP37 3 7 0.25E-12
CP24 2 4 0.24E-12
CP14 1 4 0.84E-12
RVG 1 4 13.7E6
VO 2 9 5.0E-3
Q45 10 69 57 QPC
Q46 11 60 58 QNC
Q47 56 56 8 QPC
Q48 69 69 56 QPC
Q49 60 60 59 QNC
Q50 59 59 5 QNC
RI1 8 57 1465.0
RI2 58 5 1465.0
D1 70 0 DD1
D2 71 0 DD1
IN1 0 70 1.068E-4
IN2 0 71 1.068E-4
GN1 2 4 70 71 2.0E-2
IQQ 8 5 2.0E-3
IGP 8 4 27.0E-6
Q5 16 12 14 QAP
C2 8 23 0.2E-12
I1 69 60 500.0E-6
I2 12 5 250.0E-6
R41 26 27 3.0E3
Q34 8 52 54 QN2 2
C1 0 12 3.14E-12
Q35 5 53 55 QP2 2
Q36 51 51 53 QN1
Q37 51 51 52 QP1
R53 6 54 10.0
Q3 5 9 10 QAP
R54 55 6 10.0
F5 8 23 VF5 1.0
VF5 8 22 0
Q16 8 23 26 QAN
Q14 22 1 24 QAN
Q15 23 26 24 QAN
R55 43 50 100.0
R56 42 45 100.0
C3 5 29 0.88E-12
Q41 6 45 49 QP1
Q42 43 43 44 QP1
Q4 12 3 10 QAP
F4 7 5 VF4 1.0
VF4 21 5 0
I5 13 5 250.0E-6
I9 8 30 200.0E-6
I10 8 34 100.0E-6
R45 4 36 50.0
I11 29 5 100.0E-6
F1 8 18 VF1 1.0
VF1 8 15 0
I14 8 35 500.0E-6
F3 17 5 VF3 1.0
VF3 16 5 0
I15 37 5 500.0E-6
F2 8 19 VF2 1.0
VF2 8 17 0
Q6 15 14 3 QNB
F6 43 5 VF6 4.0
VF6 38 5 0
F7 8 42 VF7 4.0
VF7 8 41 0
Q10 21 20 18 QIP
Q7 15 12 13 QAN
Q11 5 4 19 QIP
Q17 28 4 30 QAP
I6 8 14 250.0E-6
Q12 5 4 18 QIP
Q18 29 27 30 QAP
Q13 7 20 19 QIP
Q19 5 29 28 QAP
Q20 5 29 32 QAP
Q21 33 33 34 QAP
Q38 8 49 52 QN1
Q22 5 32 20 QAP
F8 48 5 VF8 1.0
VF8 47 5 0
I7 24 5 200.0E-6
Q8 16 13 3 QPB
I8 26 5 100.0E-6
Q43 42 42 44 QN1
F9 8 49 VF9 1.0
VF9 8 46 0
Q24 33 33 32 QAN
Q25 8 34 20 QAN
I3 8 12 250.0E-6
Q9 35 35 36 QAN
Q39 6 50 48 QN1
Q23 40 35 7 QAN
Q40 5 48 53 QP1
Q1 8 9 11 QAN
Q29 37 37 36 QAP
R49 38 39 37.0
R50 39 47 37.0
R51 40 41 37.0
R52 40 46 37.0
R43 27 20 1.0E3
Q30 39 37 7 QAP
R44 4 27 1.0E3
C4  5 44  0.64E-12
I13 27 5 355.0E-6
Q2 12 3 11 QAN
.MODEL DD1 D IS=1.0E-16
.MODEL QAN NPN
+ IS =0.166F    BF =3.239E+02  NF =1.000E+00  VAF=84.6
+ IKF=2.462E-02 ISE=2.956E-17  NE =1.197E+00  BR =3.719E+01
+ NR =1.000E+00 VAR=1.696E+00  IKR=3.964E-02  ISC=1.835E-19
+ NC =1.700E+00 RB =68         IRB=0.000E+00  RBM=15.1
+ RC =2.645E+01 CJE=1.632E-13  VJE=7.973E-01
+ MJE=4.950E-01 TF =1.948E-11  XTF=1.873E+01  VTF=2.825E+00
+ ITF=5.955E-02 PTF=0.000E+00  CJC=1.720E-13  VJC=8.046E-01
+ MJC=4.931E-01 XCJC=171M      TR =4.212E-10  CJS=629F
+ MJS=0         KF =100F       AF =1.000E+00
+ FC =9.765E-01
.MODEL QIP PNP
+ IS =0.166F    BF =3.239E+02 NF =1.000E+00 BR =3.719E+01
+ NR =1.000E+00 RB =68        IRB=0.000E+00 RBM=15.1
+ RC =2.645E+01 CJE=1.632E-13 VJE=7.973E-01
+ MJE=4.950E-01 TF =1.948E-11 XTF=1.873E+01 VTF=2.825E+00
+ ITF=5.955E-02 PTF=0.000E+00 CJC=1.720E-13 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=171M     TR =4.212E-10 CJS=629F
+ MJS=0         KF =100F      AF =1.000E+00 FC =9.765E-01
.MODEL QN1 NPN
+ IS =7.822E-16 BF =3.239E+02  NF =1.000E+00 VAF=8.457E+01
+ IKF=9.079E-02 ISE=1.090E-16  NE =1.197E+00 BR =3.960E+01
+ NR =1.000E+00 VAR=1.696E+00  IKR=1.462E-01 ISC=5.656E-19
+ NC =1.700E+00 RB =1.843E+01  IRB=0.000E+00 RBM=4.083E+00
+ RC =6.141E+00 CJE=5.858E-13  VJE=7.973E-01
+ MJE=4.950E-01 TF =1.874E-11  XTF=1.873E+01 VTF=2.825E+00
+ ITF=2.196E-01 PTF=0.000E+00  CJC=5.143E-13 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=1.709E-01 TR =1.069E-09 CJS=8.567E-13
+ VJS=5.723E-01 MJS=4.105E-01  KF =100F      AF =1.000E+00
+ FC =9.765E-01
.MODEL QN2 NPN
+ IS =1.880E-15 BF =1.810E+02 NF =1.000E+00 VAF=8.457E+01
+ IKF=6.800E-02 ISE=2.620E-16 NE =1.197E+00 BR =3.971E+01
+ NR =1.000E+00 VAR=1.696E+00 IKR=3.513E-01 ISC=1.348E-18
+ NC =1.700E+00 RB =57.7      IRB=0.000E+00 RBM=51.7
+ RC =3.738E+00 CJE=1.408E-12 VJE=7.973E-01
+ MJE=4.950E-01 TF =1.871E-11 XTF=1.873E+01 VTF=2.825E+00
+ ITF=5.278E-01 PTF=0.000E+00 CJC=1.224E-12 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=800M     TR =1.296E-09 CJS=1.496E-12
+ MJS=4.105E-01 KF =100F      AF =1.000E+00
+ FC =9.765E-01
.MODEL QAP PNP
+ IS =0.166F    BF =7.165E+01 NF =1.000E+00 VAF=3.439E+01
+ IKF=1.882E-02 ISE=6.380E-16 NE =1.366E+00 BR =1.833E+01
+ NR =1.000E+00 VAR=1.805E+00 IKR=1.321E-01 ISC=3.666E-18
+ NC =1.634E+00 RB =28.8      IRB=0.000E+00 RBM=7.6
+ RC =3.739E+01 CJE=1.588E-13 VJE=7.975E-01
+ MJE=5.000E-01 TF =3.156E-11 XTF=5.386E+00 VTF=2.713E+00
+ ITF=5.084E-02 PTF=0.000E+00 CJC=2.725E-13 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=170M     TR =7.500E-11 CJS=515F
+ MJS=0         KF =100F      AF =1.000E+00 FC =8.803E-01
.MODEL QP1 PNP
+ IS =4.744E-16 BF =7.165E+01  NF =1.000E+00 VAF=3.439E+01
+ IKF=6.940E-02 ISE=2.353E-15  NE =1.366E+00 BR =1.948E+01
+ NR =1.000E+00 VAR=1.805E+00  IKR=4.873E-01 ISC=1.322E-17
+ NC =1.634E+00 RB =7.797E+00  IRB=0.000E+00 RBM=2.052E+00
+ RC =1.037E+01 CJE=5.858E-13  VJE=7.975E-01
+ MJE=5.000E-01 TF =3.073E-11  XTF=5.386E+00 VTF=2.713E+00
+ ITF=1.875E-01 PTF=0.000E+00  CJC=8.147E-13 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=1.709E-01 TR =1.450E-10 CJS=1.364E-12
+ VJS=6.691E-01 MJS=3.950E-01  KF =100F      AF =1.000E+00
+ FC =8.803E-01
.MODEL QP2 PNP
+ IS =1.140E-15 BF =5.165E+01 NF =1.000E+00 VAF=3.439E+01
+ IKF=6.700E-02 ISE=5.655E-15 NE =1.366E+00 BR =1.953E+01
+ NR =1.000E+00 VAR=1.805E+00 IKR=1.171E+00 ISC=3.173E-17
+ NC =1.634E+00 RB =53.2      IRB=0.000E+00 RBM=50.9
+ RC =6.213E+00 CJE=1.408E-12 VJE=7.975E-01
+ MJE=5.000E-01 TF =3.070E-11 XTF=5.386E+00 VTF=2.713E+00
+ ITF=4.506E-01 PTF=0.000E+00 CJC=1.939E-12 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=900M     TR =1.850E-10 CJS=2.351E-12
+ MJS=3.950E-01 KF =100F      AF =1.000E+00
+ FC =8.803E-01
.MODEL QPB PNP
+ IS =4.744E-16 BF =7.165E+01  NF =1.000E+00 VAF=3.439E+01
+ IKF=7.940E-03 ISE=2.353E-15  NE =1.366E+00 BR =1.948E+01
+ NR =1.000E+00 VAR=1.805E+00  IKR=4.873E-01 ISC=1.322E-17
+ NC =1.634E+00 RB =7.797E+00  IRB=0.000E+00 RBM=2.052E+00
+ RC =1.037E+01 CJE=5.858E-13  VJE=7.975E-01
+ MJE=5.000E-01 TF =3.073E-11  XTF=5.386E+00 VTF=2.713E+00
+ ITF=1.875E-01 PTF=0.000E+00  CJC=8.147E-13 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=1.709E-01 TR =1.450E-10 CJS=1.364E-12
+ VJS=6.691E-01 MJS=3.950E-01  KF =100F      AF =1.000E+00
+ FC =8.803E-01
.MODEL QNB NPN
+ IS =7.822E-16 BF =1.039E+02  NF =1.000E+00 VAF=8.457E+01
+ IKF=8.079E-03 ISE=1.090E-16  NE =1.197E+00 BR =3.960E+01
+ NR =1.000E+00 VAR=1.696E+00  IKR=1.462E-01 ISC=5.656E-19
+ NC =1.700E+00 RB =1.843E+01  IRB=0.000E+00 RBM=4.083E+00
+ RC =6.141E+00 CJE=5.858E-13  VJE=7.973E-01
+ MJE=4.950E-01 TF =1.874E-11  XTF=1.873E+01 VTF=2.825E+00
+ ITF=2.196E-01 PTF=0.000E+00  CJC=5.143E-13 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=1.709E-01 TR =1.069E-09 CJS=8.567E-13
+ VJS=5.723E-01 MJS=4.105E-01  KF =100F      AF =1.000E+00
+ FC =9.765E-01
.MODEL QPC PNP
+ IS =4.744E-16 BF =1.000E+02  NF =1.000E+00 VAF=3.439E+01
+ IKF=7.940E-03 ISE=2.353E-15  NE =1.366E+00 BR =1.948E+01
+ NR =1.000E+00 VAR=1.805E+00  IKR=4.873E-01 ISC=1.322E-17
+ NC =1.634E+00 RB =7.797E+00  IRB=0.000E+00 RBM=2.052E+00
+ RC =1.037E+01 CJE=5.858E-13  VJE=7.975E-01
+ MJE=5.000E-01 TF =3.073E-11  XTF=5.386E+00 VTF=2.713E+00
+ ITF=1.875E-01 PTF=0.000E+00  CJC=8.147E-13 VJC=7.130E-01
+ MJC=4.200E-01 XCJC=1.709E-01 TR =1.450E-10 CJS=1.364E-12
+ VJS=6.691E-01 MJS=3.950E-01  KF =100F      AF =1.000E+00
+ FC =8.803E-01
.MODEL QNC NPN
+ IS =7.822E-16 BF =1.000E+02  NF =1.000E+00 VAF=8.457E+01
+ IKF=8.079E-03 ISE=1.090E-16  NE =1.197E+00 BR =3.960E+01
+ NR =1.000E+00 VAR=1.696E+00  IKR=1.462E-01 ISC=5.656E-19
+ NC =1.700E+00 RB =1.843E+01  IRB=0.000E+00 RBM=4.083E+00
+ RC =6.141E+00 CJE=5.858E-13  VJE=7.973E-01
+ MJE=4.950E-01 TF =1.874E-11  XTF=1.873E+01 VTF=2.825E+00
+ ITF=2.196E-01 PTF=0.000E+00  CJC=5.143E-13 VJC=8.046E-01
+ MJC=4.931E-01 XCJC=1.709E-01 TR =1.069E-09 CJS=8.567E-13
+ VJS=5.723E-01 MJS=4.105E-01  KF =100F      AF =1.000E+00
+ FC =9.765E-01
.ENDS

