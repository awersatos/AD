*  
* Diode Model Produced by Altium Ltd  
* Date:  4-May-2004 
*  
* Manufacturer: Renesas  
* Component Name: HDSP-503B  
*  
* Parameters derived from information available in data sheet.  
*
*                 anode-e
*                 |  anode-d
*                 |  |  common-cathode
*                 |  |  |  anode-c
*                 |  |  |  |  anode-DP
*                 |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  |  |  anode-f
*                 |  |  |  |  |  |  |  |  |  anode-g
*                 |  |  |  |  |  |  |  |  |  |  
.SUBCKT HDSP_503B 1  2  3  4  5  6  7  8  9  10

DA1   7  3  dHDSP_503B
DB1   6  3  dHDSP_503B
DC1   4  3  dHDSP_503B
DD1   2  3  dHDSP_503B
DE1   1  3  dHDSP_503B
DF1   9  3  dHDSP_503B
DG1  10  3  dHDSP_503B
DDP1  5  3  dHDSP_503B

DA2   7  8  dHDSP_503B
DB2   6  8  dHDSP_503B
DC2   4  8  dHDSP_503B
DD2   2  8  dHDSP_503B
DE2   1  8  dHDSP_503B
DF2   9  8  dHDSP_503B
DG2  10  8  dHDSP_503B
DDP2  5  8  dHDSP_503B

.MODEL dHDSP_503B D
+ (  
+    IS = 2.15137703E-17 
+    N  = 4.02940472 
+    RS = 16.32357710 
+    BV = 4.50000000 
+    IBV = 100u 
+ )  

.ENDS HDSP_503B