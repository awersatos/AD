*DPDT Relay Subcircuit Parameters
*PULLIN     = Pull in voltage
*DROPOFF    = Drop off voltage
*CONTACT    = Contact resistance
*RESISTANCE = Coil resistance
*INDUCTANCE = Coil Inductance 
* jjt 15/6/2002: extended existing SPDT model to DPDT.
*
*Generic DPDT Relay
*Connections:     COM1
*                 | NC1
*                 | | NO1
*                 | | | T1
*                 | | | | T2
*                 | | | | | COM2
*                 | | | | | |  NC2
*                 | | | | | |  |  NO2
*                 | | | | | |  |  |
*                 | | | | | |  |  |
.SUBCKT DPDTRELAY 1 2 3 4 5 11 12 13
+ PARAMS: PULLIN=4 DROPOFF=0.1 CONTACT=1m RESISTANCE=500 INDUCTANCE=10m
L1 4 6 {(INDUCTANCE/2)}
L2 5 7 {(INDUCTANCE/2)}
R1 6 7 {RESISTANCE}
*
BNO1 8 0 V={PULLIN}-abs(v(6,7))
SW1 2 1 8 0 SWNC ON
BNC1 9 0 V=abs(v(6,7))
SW2 3 1 9 0 SWNO OFF
*
BNO2 15 0 V={PULLIN}-abs(v(6,7))
SW3 12 11 15 0 SWNC ON
BNC2 16 0 V=abs(v(6,7))
SW4 13 11 16 0 SWNO OFF
*
.MODEL SWNC SW(VT={DROPOFF} RON={CONTACT} )
.MODEL SWNO SW(VT={(PULLIN*0.98)} RON={CONTACT} )
.ENDS DPDTRELAY