-------------------------------------------------------------------------------
-- This is an automatically generated file. 
-- Note some spartan3/6 work-arounds added manually.
-------------------------------------------------------------------------------
--   ____  ____
--  /   /\/   /
-- /___/  \  /   Vendor: Xilinx
-- \   \   \/    Version: 4.0
--  \   \        Filename: $RCSfile: dds_compiler_v4_0_eff_lut.vhd,v $
--  /   /        Date Last Modified: $Date: 2009/12/04 11:46:31 $
-- /___/   /\    Date Created: 2009
-- \   \  /  \
--  \___\/\___\
--
-- Device  : All
-- Library : dds_compiler_v4_0
-- Purpose : LUT to calculate ((x-0.5)*pi)^2
-------------------------------------------------------------------------------
--  (c) Copyright 2009 Xilinx, Inc. All rights reserved.
--
--  This file contains confidential and proprietary information
--  of Xilinx, Inc. and is protected under U.S. and
--  international copyright and other intellectual property
--  laws.
--
--  DISCLAIMER
--  This disclaimer is not a license and does not grant any
--  rights to the materials distributed herewith. Except as
--  otherwise provided in a valid license issued to you by
--  Xilinx, and to the maximum extent permitted by applicable
--  law: (1) THESE MATERIALS ARE MADE AVAILABLE "AS IS" AND
--  WITH ALL FAULTS, AND XILINX HEREBY DISCLAIMS ALL WARRANTIES
--  AND CONDITIONS, EXPRESS, IMPLIED, OR STATUTORY, INCLUDING
--  BUT NOT LIMITED TO WARRANTIES OF MERCHANTABILITY, NON-
--  INFRINGEMENT, OR FITNESS FOR ANY PARTICULAR PURPOSE; and
--  (2) Xilinx shall not be liable (whether in contract or tort,
--  including negligence, or under any other theory of
--  liability) for any loss or damage of any kind or nature
--  related to, arising under or in connection with these
--  materials, including for any direct, or any indirect,
--  special, incidental, or consequential loss or damage
--  (including loss of data, profits, goodwill, or any type of
--  loss or damage suffered as a result of any action brought
--  by a third party) even if such damage or loss was
--  reasonably foreseeable or Xilinx had been advised of the
--  possibility of the same.
--
--  CRITICAL APPLICATIONS
--  Xilinx products are not designed or intended to be fail-
--  safe, or for use in any application requiring fail-safe
--  performance, such as life-support or safety devices or
--  systems, Class III medical devices, nuclear facilities,
--  applications related to the deployment of airbags, or any
--  other applications that could lead to death, personal
--  injury, or severe property or environmental damage
--  (individually and collectively, "Critical
--  Applications"). Customer assumes the sole risk and
--  liability of any use of Xilinx products in Critical
--  Applications, subject only to applicable laws and
--  regulations governing limitations on product liability.
--
--  THIS COPYRIGHT NOTICE AND DISCLAIMER MUST BE RETAINED AS
--  PART OF THIS FILE AT ALL TIMES.
-------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library xilinxcorelib;
use xilinxcorelib.bip_utils_pkg_v2_0.all;

library xilinxcorelib;
use xilinxcorelib.xbip_pipe_v2_0_xst_comp.all;

library xilinxcorelib;
use xilinxcorelib.xbip_bram18k_v2_1_xst_comp.all;
use xilinxcorelib.bip_bram18k_pkg_v2_1.all;
use xilinxcorelib.bip_bram18k_v2_1_sim_pkg.all;

entity dds_compiler_v4_0_eff_lut is
 generic (
    C_XDEVICEFAMILY : string  := "virtex4";
    C_LATENCY       : integer := -1;
    C_MODEL_TYPE    : integer := 0          -- 0 = synth, 1 = RTL
    );
  port (
    CLK             : in  std_logic := '1';
    CE              : in  std_logic := '1';
    SCLR            : in  std_logic := '0';
    A               : in  std_logic_vector(9 downto 0)  := (others => '0');
    D               : out std_logic_vector(17 downto 0) := (others => '0')
    );
  end dds_compiler_v4_0_eff_lut;

  architecture rtl of dds_compiler_v4_0_eff_lut is

  constant ci_data_table : t_BRAM18k_10_18_init_val := (
    "000000010011101111",  -- (p-0.5)^2*pi^2(0.00)=2.467401e+00
    "000000010011101010",  -- (p-0.5)^2*pi^2(0.00)=2.457772e+00
    "000000010011100101",  -- (p-0.5)^2*pi^2(0.00)=2.448162e+00
    "000000010011100001",  -- (p-0.5)^2*pi^2(0.00)=2.438571e+00
    "000000010011011100",  -- (p-0.5)^2*pi^2(0.00)=2.428999e+00
    "000000010011010111",  -- (p-0.5)^2*pi^2(0.00)=2.419445e+00
    "000000010011010010",  -- (p-0.5)^2*pi^2(0.01)=2.409910e+00
    "000000010011001101",  -- (p-0.5)^2*pi^2(0.01)=2.400394e+00
    "000000010011001000",  -- (p-0.5)^2*pi^2(0.01)=2.390897e+00
    "000000010011000011",  -- (p-0.5)^2*pi^2(0.01)=2.381419e+00
    "000000010010111110",  -- (p-0.5)^2*pi^2(0.01)=2.371959e+00
    "000000010010111010",  -- (p-0.5)^2*pi^2(0.01)=2.362519e+00
    "000000010010110101",  -- (p-0.5)^2*pi^2(0.01)=2.353097e+00
    "000000010010110000",  -- (p-0.5)^2*pi^2(0.01)=2.343694e+00
    "000000010010101011",  -- (p-0.5)^2*pi^2(0.01)=2.334310e+00
    "000000010010100110",  -- (p-0.5)^2*pi^2(0.01)=2.324945e+00
    "000000010010100010",  -- (p-0.5)^2*pi^2(0.02)=2.315598e+00
    "000000010010011101",  -- (p-0.5)^2*pi^2(0.02)=2.306270e+00
    "000000010010011000",  -- (p-0.5)^2*pi^2(0.02)=2.296962e+00
    "000000010010010011",  -- (p-0.5)^2*pi^2(0.02)=2.287672e+00
    "000000010010001111",  -- (p-0.5)^2*pi^2(0.02)=2.278400e+00
    "000000010010001010",  -- (p-0.5)^2*pi^2(0.02)=2.269148e+00
    "000000010010000101",  -- (p-0.5)^2*pi^2(0.02)=2.259914e+00
    "000000010010000000",  -- (p-0.5)^2*pi^2(0.02)=2.250700e+00
    "000000010001111100",  -- (p-0.5)^2*pi^2(0.02)=2.241504e+00
    "000000010001110111",  -- (p-0.5)^2*pi^2(0.02)=2.232327e+00
    "000000010001110010",  -- (p-0.5)^2*pi^2(0.03)=2.223168e+00
    "000000010001101110",  -- (p-0.5)^2*pi^2(0.03)=2.214029e+00
    "000000010001101001",  -- (p-0.5)^2*pi^2(0.03)=2.204908e+00
    "000000010001100100",  -- (p-0.5)^2*pi^2(0.03)=2.195807e+00
    "000000010001100000",  -- (p-0.5)^2*pi^2(0.03)=2.186724e+00
    "000000010001011011",  -- (p-0.5)^2*pi^2(0.03)=2.177660e+00
    "000000010001010110",  -- (p-0.5)^2*pi^2(0.03)=2.168614e+00
    "000000010001010010",  -- (p-0.5)^2*pi^2(0.03)=2.159588e+00
    "000000010001001101",  -- (p-0.5)^2*pi^2(0.03)=2.150580e+00
    "000000010001001000",  -- (p-0.5)^2*pi^2(0.03)=2.141591e+00
    "000000010001000100",  -- (p-0.5)^2*pi^2(0.04)=2.132621e+00
    "000000010000111111",  -- (p-0.5)^2*pi^2(0.04)=2.123670e+00
    "000000010000111011",  -- (p-0.5)^2*pi^2(0.04)=2.114738e+00
    "000000010000110110",  -- (p-0.5)^2*pi^2(0.04)=2.105824e+00
    "000000010000110010",  -- (p-0.5)^2*pi^2(0.04)=2.096929e+00
    "000000010000101101",  -- (p-0.5)^2*pi^2(0.04)=2.088054e+00
    "000000010000101001",  -- (p-0.5)^2*pi^2(0.04)=2.079197e+00
    "000000010000100100",  -- (p-0.5)^2*pi^2(0.04)=2.070358e+00
    "000000010000100000",  -- (p-0.5)^2*pi^2(0.04)=2.061539e+00
    "000000010000011011",  -- (p-0.5)^2*pi^2(0.04)=2.052738e+00
    "000000010000010111",  -- (p-0.5)^2*pi^2(0.04)=2.043957e+00
    "000000010000010010",  -- (p-0.5)^2*pi^2(0.05)=2.035194e+00
    "000000010000001110",  -- (p-0.5)^2*pi^2(0.05)=2.026450e+00
    "000000010000001001",  -- (p-0.5)^2*pi^2(0.05)=2.017724e+00
    "000000010000000101",  -- (p-0.5)^2*pi^2(0.05)=2.009018e+00
    "000000010000000000",  -- (p-0.5)^2*pi^2(0.05)=2.000330e+00
    "000000001111111100",  -- (p-0.5)^2*pi^2(0.05)=1.991661e+00
    "000000001111110111",  -- (p-0.5)^2*pi^2(0.05)=1.983011e+00
    "000000001111110011",  -- (p-0.5)^2*pi^2(0.05)=1.974380e+00
    "000000001111101110",  -- (p-0.5)^2*pi^2(0.05)=1.965768e+00
    "000000001111101010",  -- (p-0.5)^2*pi^2(0.05)=1.957174e+00
    "000000001111100110",  -- (p-0.5)^2*pi^2(0.06)=1.948600e+00
    "000000001111100001",  -- (p-0.5)^2*pi^2(0.06)=1.940044e+00
    "000000001111011101",  -- (p-0.5)^2*pi^2(0.06)=1.931507e+00
    "000000001111011001",  -- (p-0.5)^2*pi^2(0.06)=1.922989e+00
    "000000001111010100",  -- (p-0.5)^2*pi^2(0.06)=1.914489e+00
    "000000001111010000",  -- (p-0.5)^2*pi^2(0.06)=1.906009e+00
    "000000001111001100",  -- (p-0.5)^2*pi^2(0.06)=1.897547e+00
    "000000001111000111",  -- (p-0.5)^2*pi^2(0.06)=1.889104e+00
    "000000001111000011",  -- (p-0.5)^2*pi^2(0.06)=1.880680e+00
    "000000001110111111",  -- (p-0.5)^2*pi^2(0.06)=1.872275e+00
    "000000001110111010",  -- (p-0.5)^2*pi^2(0.07)=1.863888e+00
    "000000001110110110",  -- (p-0.5)^2*pi^2(0.07)=1.855521e+00
    "000000001110110010",  -- (p-0.5)^2*pi^2(0.07)=1.847172e+00
    "000000001110101101",  -- (p-0.5)^2*pi^2(0.07)=1.838842e+00
    "000000001110101001",  -- (p-0.5)^2*pi^2(0.07)=1.830531e+00
    "000000001110100101",  -- (p-0.5)^2*pi^2(0.07)=1.822238e+00
    "000000001110100001",  -- (p-0.5)^2*pi^2(0.07)=1.813965e+00
    "000000001110011101",  -- (p-0.5)^2*pi^2(0.07)=1.805710e+00
    "000000001110011000",  -- (p-0.5)^2*pi^2(0.07)=1.797474e+00
    "000000001110010100",  -- (p-0.5)^2*pi^2(0.07)=1.789257e+00
    "000000001110010000",  -- (p-0.5)^2*pi^2(0.08)=1.781059e+00
    "000000001110001100",  -- (p-0.5)^2*pi^2(0.08)=1.772880e+00
    "000000001110001000",  -- (p-0.5)^2*pi^2(0.08)=1.764719e+00
    "000000001110000011",  -- (p-0.5)^2*pi^2(0.08)=1.756578e+00
    "000000001101111111",  -- (p-0.5)^2*pi^2(0.08)=1.748455e+00
    "000000001101111011",  -- (p-0.5)^2*pi^2(0.08)=1.740351e+00
    "000000001101110111",  -- (p-0.5)^2*pi^2(0.08)=1.732265e+00
    "000000001101110011",  -- (p-0.5)^2*pi^2(0.08)=1.724199e+00
    "000000001101101111",  -- (p-0.5)^2*pi^2(0.08)=1.716151e+00
    "000000001101101011",  -- (p-0.5)^2*pi^2(0.08)=1.708123e+00
    "000000001101100110",  -- (p-0.5)^2*pi^2(0.08)=1.700113e+00
    "000000001101100010",  -- (p-0.5)^2*pi^2(0.09)=1.692122e+00
    "000000001101011110",  -- (p-0.5)^2*pi^2(0.09)=1.684149e+00
    "000000001101011010",  -- (p-0.5)^2*pi^2(0.09)=1.676196e+00
    "000000001101010110",  -- (p-0.5)^2*pi^2(0.09)=1.668261e+00
    "000000001101010010",  -- (p-0.5)^2*pi^2(0.09)=1.660345e+00
    "000000001101001110",  -- (p-0.5)^2*pi^2(0.09)=1.652448e+00
    "000000001101001010",  -- (p-0.5)^2*pi^2(0.09)=1.644570e+00
    "000000001101000110",  -- (p-0.5)^2*pi^2(0.09)=1.636711e+00
    "000000001101000010",  -- (p-0.5)^2*pi^2(0.09)=1.628870e+00
    "000000001100111110",  -- (p-0.5)^2*pi^2(0.09)=1.621049e+00
    "000000001100111010",  -- (p-0.5)^2*pi^2(0.10)=1.613246e+00
    "000000001100110110",  -- (p-0.5)^2*pi^2(0.10)=1.605462e+00
    "000000001100110010",  -- (p-0.5)^2*pi^2(0.10)=1.597696e+00
    "000000001100101110",  -- (p-0.5)^2*pi^2(0.10)=1.589950e+00
    "000000001100101010",  -- (p-0.5)^2*pi^2(0.10)=1.582222e+00
    "000000001100100110",  -- (p-0.5)^2*pi^2(0.10)=1.574514e+00
    "000000001100100010",  -- (p-0.5)^2*pi^2(0.10)=1.566824e+00
    "000000001100011110",  -- (p-0.5)^2*pi^2(0.10)=1.559153e+00
    "000000001100011010",  -- (p-0.5)^2*pi^2(0.10)=1.551500e+00
    "000000001100010110",  -- (p-0.5)^2*pi^2(0.10)=1.543867e+00
    "000000001100010011",  -- (p-0.5)^2*pi^2(0.11)=1.536252e+00
    "000000001100001111",  -- (p-0.5)^2*pi^2(0.11)=1.528657e+00
    "000000001100001011",  -- (p-0.5)^2*pi^2(0.11)=1.521080e+00
    "000000001100000111",  -- (p-0.5)^2*pi^2(0.11)=1.513521e+00
    "000000001100000011",  -- (p-0.5)^2*pi^2(0.11)=1.505982e+00
    "000000001011111111",  -- (p-0.5)^2*pi^2(0.11)=1.498462e+00
    "000000001011111011",  -- (p-0.5)^2*pi^2(0.11)=1.490960e+00
    "000000001011111000",  -- (p-0.5)^2*pi^2(0.11)=1.483477e+00
    "000000001011110100",  -- (p-0.5)^2*pi^2(0.11)=1.476013e+00
    "000000001011110000",  -- (p-0.5)^2*pi^2(0.11)=1.468568e+00
    "000000001011101100",  -- (p-0.5)^2*pi^2(0.12)=1.461141e+00
    "000000001011101000",  -- (p-0.5)^2*pi^2(0.12)=1.453734e+00
    "000000001011100101",  -- (p-0.5)^2*pi^2(0.12)=1.446345e+00
    "000000001011100001",  -- (p-0.5)^2*pi^2(0.12)=1.438975e+00
    "000000001011011101",  -- (p-0.5)^2*pi^2(0.12)=1.431624e+00
    "000000001011011001",  -- (p-0.5)^2*pi^2(0.12)=1.424292e+00
    "000000001011010101",  -- (p-0.5)^2*pi^2(0.12)=1.416979e+00
    "000000001011010010",  -- (p-0.5)^2*pi^2(0.12)=1.409684e+00
    "000000001011001110",  -- (p-0.5)^2*pi^2(0.12)=1.402408e+00
    "000000001011001010",  -- (p-0.5)^2*pi^2(0.12)=1.395151e+00
    "000000001011000111",  -- (p-0.5)^2*pi^2(0.12)=1.387913e+00
    "000000001011000011",  -- (p-0.5)^2*pi^2(0.13)=1.380694e+00
    "000000001010111111",  -- (p-0.5)^2*pi^2(0.13)=1.373493e+00
    "000000001010111100",  -- (p-0.5)^2*pi^2(0.13)=1.366312e+00
    "000000001010111000",  -- (p-0.5)^2*pi^2(0.13)=1.359149e+00
    "000000001010110100",  -- (p-0.5)^2*pi^2(0.13)=1.352005e+00
    "000000001010110001",  -- (p-0.5)^2*pi^2(0.13)=1.344880e+00
    "000000001010101101",  -- (p-0.5)^2*pi^2(0.13)=1.337773e+00
    "000000001010101001",  -- (p-0.5)^2*pi^2(0.13)=1.330686e+00
    "000000001010100110",  -- (p-0.5)^2*pi^2(0.13)=1.323617e+00
    "000000001010100010",  -- (p-0.5)^2*pi^2(0.13)=1.316567e+00
    "000000001010011110",  -- (p-0.5)^2*pi^2(0.14)=1.309536e+00
    "000000001010011011",  -- (p-0.5)^2*pi^2(0.14)=1.302524e+00
    "000000001010010111",  -- (p-0.5)^2*pi^2(0.14)=1.295531e+00
    "000000001010010100",  -- (p-0.5)^2*pi^2(0.14)=1.288556e+00
    "000000001010010000",  -- (p-0.5)^2*pi^2(0.14)=1.281600e+00
    "000000001010001101",  -- (p-0.5)^2*pi^2(0.14)=1.274663e+00
    "000000001010001001",  -- (p-0.5)^2*pi^2(0.14)=1.267745e+00
    "000000001010000110",  -- (p-0.5)^2*pi^2(0.14)=1.260846e+00
    "000000001010000010",  -- (p-0.5)^2*pi^2(0.14)=1.253965e+00
    "000000001001111111",  -- (p-0.5)^2*pi^2(0.14)=1.247104e+00
    "000000001001111011",  -- (p-0.5)^2*pi^2(0.15)=1.240261e+00
    "000000001001111000",  -- (p-0.5)^2*pi^2(0.15)=1.233437e+00
    "000000001001110100",  -- (p-0.5)^2*pi^2(0.15)=1.226632e+00
    "000000001001110001",  -- (p-0.5)^2*pi^2(0.15)=1.219846e+00
    "000000001001101101",  -- (p-0.5)^2*pi^2(0.15)=1.213078e+00
    "000000001001101010",  -- (p-0.5)^2*pi^2(0.15)=1.206329e+00
    "000000001001100110",  -- (p-0.5)^2*pi^2(0.15)=1.199599e+00
    "000000001001100011",  -- (p-0.5)^2*pi^2(0.15)=1.192888e+00
    "000000001001011111",  -- (p-0.5)^2*pi^2(0.15)=1.186196e+00
    "000000001001011100",  -- (p-0.5)^2*pi^2(0.15)=1.179523e+00
    "000000001001011001",  -- (p-0.5)^2*pi^2(0.16)=1.172868e+00
    "000000001001010101",  -- (p-0.5)^2*pi^2(0.16)=1.166233e+00
    "000000001001010010",  -- (p-0.5)^2*pi^2(0.16)=1.159616e+00
    "000000001001001110",  -- (p-0.5)^2*pi^2(0.16)=1.153018e+00
    "000000001001001011",  -- (p-0.5)^2*pi^2(0.16)=1.146438e+00
    "000000001001001000",  -- (p-0.5)^2*pi^2(0.16)=1.139878e+00
    "000000001001000100",  -- (p-0.5)^2*pi^2(0.16)=1.133336e+00
    "000000001001000001",  -- (p-0.5)^2*pi^2(0.16)=1.126813e+00
    "000000001000111110",  -- (p-0.5)^2*pi^2(0.16)=1.120310e+00
    "000000001000111010",  -- (p-0.5)^2*pi^2(0.16)=1.113824e+00
    "000000001000110111",  -- (p-0.5)^2*pi^2(0.17)=1.107358e+00
    "000000001000110100",  -- (p-0.5)^2*pi^2(0.17)=1.100911e+00
    "000000001000110000",  -- (p-0.5)^2*pi^2(0.17)=1.094482e+00
    "000000001000101101",  -- (p-0.5)^2*pi^2(0.17)=1.088072e+00
    "000000001000101010",  -- (p-0.5)^2*pi^2(0.17)=1.081681e+00
    "000000001000100111",  -- (p-0.5)^2*pi^2(0.17)=1.075309e+00
    "000000001000100011",  -- (p-0.5)^2*pi^2(0.17)=1.068956e+00
    "000000001000100000",  -- (p-0.5)^2*pi^2(0.17)=1.062621e+00
    "000000001000011101",  -- (p-0.5)^2*pi^2(0.17)=1.056305e+00
    "000000001000011010",  -- (p-0.5)^2*pi^2(0.17)=1.050008e+00
    "000000001000010110",  -- (p-0.5)^2*pi^2(0.17)=1.043730e+00
    "000000001000010011",  -- (p-0.5)^2*pi^2(0.18)=1.037471e+00
    "000000001000010000",  -- (p-0.5)^2*pi^2(0.18)=1.031231e+00
    "000000001000001101",  -- (p-0.5)^2*pi^2(0.18)=1.025009e+00
    "000000001000001010",  -- (p-0.5)^2*pi^2(0.18)=1.018806e+00
    "000000001000000110",  -- (p-0.5)^2*pi^2(0.18)=1.012622e+00
    "000000001000000011",  -- (p-0.5)^2*pi^2(0.18)=1.006457e+00
    "000000001000000000",  -- (p-0.5)^2*pi^2(0.18)=1.000311e+00
    "000000000111111101",  -- (p-0.5)^2*pi^2(0.18)=9.941835e-01
    "000000000111111010",  -- (p-0.5)^2*pi^2(0.18)=9.880749e-01
    "000000000111110111",  -- (p-0.5)^2*pi^2(0.18)=9.819851e-01
    "000000000111110100",  -- (p-0.5)^2*pi^2(0.19)=9.759141e-01
    "000000000111110001",  -- (p-0.5)^2*pi^2(0.19)=9.698619e-01
    "000000000111101101",  -- (p-0.5)^2*pi^2(0.19)=9.638286e-01
    "000000000111101010",  -- (p-0.5)^2*pi^2(0.19)=9.578140e-01
    "000000000111100111",  -- (p-0.5)^2*pi^2(0.19)=9.518183e-01
    "000000000111100100",  -- (p-0.5)^2*pi^2(0.19)=9.458415e-01
    "000000000111100001",  -- (p-0.5)^2*pi^2(0.19)=9.398834e-01
    "000000000111011110",  -- (p-0.5)^2*pi^2(0.19)=9.339442e-01
    "000000000111011011",  -- (p-0.5)^2*pi^2(0.19)=9.280238e-01
    "000000000111011000",  -- (p-0.5)^2*pi^2(0.19)=9.221223e-01
    "000000000111010101",  -- (p-0.5)^2*pi^2(0.20)=9.162395e-01
    "000000000111010010",  -- (p-0.5)^2*pi^2(0.20)=9.103756e-01
    "000000000111001111",  -- (p-0.5)^2*pi^2(0.20)=9.045305e-01
    "000000000111001100",  -- (p-0.5)^2*pi^2(0.20)=8.987042e-01
    "000000000111001001",  -- (p-0.5)^2*pi^2(0.20)=8.928968e-01
    "000000000111000110",  -- (p-0.5)^2*pi^2(0.20)=8.871082e-01
    "000000000111000011",  -- (p-0.5)^2*pi^2(0.20)=8.813384e-01
    "000000000111000000",  -- (p-0.5)^2*pi^2(0.20)=8.755874e-01
    "000000000110111101",  -- (p-0.5)^2*pi^2(0.20)=8.698553e-01
    "000000000110111010",  -- (p-0.5)^2*pi^2(0.20)=8.641420e-01
    "000000000110111000",  -- (p-0.5)^2*pi^2(0.21)=8.584475e-01
    "000000000110110101",  -- (p-0.5)^2*pi^2(0.21)=8.527718e-01
    "000000000110110010",  -- (p-0.5)^2*pi^2(0.21)=8.471149e-01
    "000000000110101111",  -- (p-0.5)^2*pi^2(0.21)=8.414769e-01
    "000000000110101100",  -- (p-0.5)^2*pi^2(0.21)=8.358577e-01
    "000000000110101001",  -- (p-0.5)^2*pi^2(0.21)=8.302574e-01
    "000000000110100110",  -- (p-0.5)^2*pi^2(0.21)=8.246758e-01
    "000000000110100011",  -- (p-0.5)^2*pi^2(0.21)=8.191131e-01
    "000000000110100001",  -- (p-0.5)^2*pi^2(0.21)=8.135692e-01
    "000000000110011110",  -- (p-0.5)^2*pi^2(0.21)=8.080441e-01
    "000000000110011011",  -- (p-0.5)^2*pi^2(0.21)=8.025379e-01
    "000000000110011000",  -- (p-0.5)^2*pi^2(0.22)=7.970504e-01
    "000000000110010101",  -- (p-0.5)^2*pi^2(0.22)=7.915819e-01
    "000000000110010010",  -- (p-0.5)^2*pi^2(0.22)=7.861321e-01
    "000000000110010000",  -- (p-0.5)^2*pi^2(0.22)=7.807011e-01
    "000000000110001101",  -- (p-0.5)^2*pi^2(0.22)=7.752890e-01
    "000000000110001010",  -- (p-0.5)^2*pi^2(0.22)=7.698957e-01
    "000000000110000111",  -- (p-0.5)^2*pi^2(0.22)=7.645212e-01
    "000000000110000101",  -- (p-0.5)^2*pi^2(0.22)=7.591656e-01
    "000000000110000010",  -- (p-0.5)^2*pi^2(0.22)=7.538288e-01
    "000000000101111111",  -- (p-0.5)^2*pi^2(0.22)=7.485108e-01
    "000000000101111101",  -- (p-0.5)^2*pi^2(0.23)=7.432116e-01
    "000000000101111010",  -- (p-0.5)^2*pi^2(0.23)=7.379312e-01
    "000000000101110111",  -- (p-0.5)^2*pi^2(0.23)=7.326697e-01
    "000000000101110100",  -- (p-0.5)^2*pi^2(0.23)=7.274270e-01
    "000000000101110010",  -- (p-0.5)^2*pi^2(0.23)=7.222031e-01
    "000000000101101111",  -- (p-0.5)^2*pi^2(0.23)=7.169981e-01
    "000000000101101100",  -- (p-0.5)^2*pi^2(0.23)=7.118119e-01
    "000000000101101010",  -- (p-0.5)^2*pi^2(0.23)=7.066445e-01
    "000000000101100111",  -- (p-0.5)^2*pi^2(0.23)=7.014959e-01
    "000000000101100101",  -- (p-0.5)^2*pi^2(0.23)=6.963661e-01
    "000000000101100010",  -- (p-0.5)^2*pi^2(0.24)=6.912552e-01
    "000000000101011111",  -- (p-0.5)^2*pi^2(0.24)=6.861631e-01
    "000000000101011101",  -- (p-0.5)^2*pi^2(0.24)=6.810898e-01
    "000000000101011010",  -- (p-0.5)^2*pi^2(0.24)=6.760354e-01
    "000000000101011000",  -- (p-0.5)^2*pi^2(0.24)=6.709997e-01
    "000000000101010101",  -- (p-0.5)^2*pi^2(0.24)=6.659829e-01
    "000000000101010010",  -- (p-0.5)^2*pi^2(0.24)=6.609850e-01
    "000000000101010000",  -- (p-0.5)^2*pi^2(0.24)=6.560058e-01
    "000000000101001101",  -- (p-0.5)^2*pi^2(0.24)=6.510455e-01
    "000000000101001011",  -- (p-0.5)^2*pi^2(0.24)=6.461040e-01
    "000000000101001000",  -- (p-0.5)^2*pi^2(0.25)=6.411813e-01
    "000000000101000110",  -- (p-0.5)^2*pi^2(0.25)=6.362774e-01
    "000000000101000011",  -- (p-0.5)^2*pi^2(0.25)=6.313924e-01
    "000000000101000001",  -- (p-0.5)^2*pi^2(0.25)=6.265262e-01
    "000000000100111110",  -- (p-0.5)^2*pi^2(0.25)=6.216788e-01
    "000000000100111100",  -- (p-0.5)^2*pi^2(0.25)=6.168503e-01
    "000000000100111001",  -- (p-0.5)^2*pi^2(0.25)=6.120405e-01
    "000000000100110111",  -- (p-0.5)^2*pi^2(0.25)=6.072496e-01
    "000000000100110100",  -- (p-0.5)^2*pi^2(0.25)=6.024776e-01
    "000000000100110010",  -- (p-0.5)^2*pi^2(0.25)=5.977243e-01
    "000000000100110000",  -- (p-0.5)^2*pi^2(0.25)=5.929899e-01
    "000000000100101101",  -- (p-0.5)^2*pi^2(0.26)=5.882743e-01
    "000000000100101011",  -- (p-0.5)^2*pi^2(0.26)=5.835775e-01
    "000000000100101000",  -- (p-0.5)^2*pi^2(0.26)=5.788995e-01
    "000000000100100110",  -- (p-0.5)^2*pi^2(0.26)=5.742404e-01
    "000000000100100100",  -- (p-0.5)^2*pi^2(0.26)=5.696001e-01
    "000000000100100001",  -- (p-0.5)^2*pi^2(0.26)=5.649786e-01
    "000000000100011111",  -- (p-0.5)^2*pi^2(0.26)=5.603759e-01
    "000000000100011101",  -- (p-0.5)^2*pi^2(0.26)=5.557921e-01
    "000000000100011010",  -- (p-0.5)^2*pi^2(0.26)=5.512271e-01
    "000000000100011000",  -- (p-0.5)^2*pi^2(0.26)=5.466809e-01
    "000000000100010110",  -- (p-0.5)^2*pi^2(0.27)=5.421536e-01
    "000000000100010011",  -- (p-0.5)^2*pi^2(0.27)=5.376450e-01
    "000000000100010001",  -- (p-0.5)^2*pi^2(0.27)=5.331553e-01
    "000000000100001111",  -- (p-0.5)^2*pi^2(0.27)=5.286844e-01
    "000000000100001100",  -- (p-0.5)^2*pi^2(0.27)=5.242324e-01
    "000000000100001010",  -- (p-0.5)^2*pi^2(0.27)=5.197991e-01
    "000000000100001000",  -- (p-0.5)^2*pi^2(0.27)=5.153847e-01
    "000000000100000110",  -- (p-0.5)^2*pi^2(0.27)=5.109891e-01
    "000000000100000011",  -- (p-0.5)^2*pi^2(0.27)=5.066124e-01
    "000000000100000001",  -- (p-0.5)^2*pi^2(0.27)=5.022544e-01
    "000000000011111111",  -- (p-0.5)^2*pi^2(0.28)=4.979153e-01
    "000000000011111101",  -- (p-0.5)^2*pi^2(0.28)=4.935951e-01
    "000000000011111011",  -- (p-0.5)^2*pi^2(0.28)=4.892936e-01
    "000000000011111000",  -- (p-0.5)^2*pi^2(0.28)=4.850110e-01
    "000000000011110110",  -- (p-0.5)^2*pi^2(0.28)=4.807471e-01
    "000000000011110100",  -- (p-0.5)^2*pi^2(0.28)=4.765022e-01
    "000000000011110010",  -- (p-0.5)^2*pi^2(0.28)=4.722760e-01
    "000000000011110000",  -- (p-0.5)^2*pi^2(0.28)=4.680687e-01
    "000000000011101110",  -- (p-0.5)^2*pi^2(0.28)=4.638801e-01
    "000000000011101011",  -- (p-0.5)^2*pi^2(0.28)=4.597105e-01
    "000000000011101001",  -- (p-0.5)^2*pi^2(0.29)=4.555596e-01
    "000000000011100111",  -- (p-0.5)^2*pi^2(0.29)=4.514276e-01
    "000000000011100101",  -- (p-0.5)^2*pi^2(0.29)=4.473143e-01
    "000000000011100011",  -- (p-0.5)^2*pi^2(0.29)=4.432199e-01
    "000000000011100001",  -- (p-0.5)^2*pi^2(0.29)=4.391444e-01
    "000000000011011111",  -- (p-0.5)^2*pi^2(0.29)=4.350876e-01
    "000000000011011101",  -- (p-0.5)^2*pi^2(0.29)=4.310497e-01
    "000000000011011011",  -- (p-0.5)^2*pi^2(0.29)=4.270306e-01
    "000000000011011001",  -- (p-0.5)^2*pi^2(0.29)=4.230304e-01
    "000000000011010111",  -- (p-0.5)^2*pi^2(0.29)=4.190489e-01
    "000000000011010101",  -- (p-0.5)^2*pi^2(0.29)=4.150863e-01
    "000000000011010011",  -- (p-0.5)^2*pi^2(0.30)=4.111425e-01
    "000000000011010000",  -- (p-0.5)^2*pi^2(0.30)=4.072176e-01
    "000000000011001110",  -- (p-0.5)^2*pi^2(0.30)=4.033114e-01
    "000000000011001101",  -- (p-0.5)^2*pi^2(0.30)=3.994241e-01
    "000000000011001011",  -- (p-0.5)^2*pi^2(0.30)=3.955556e-01
    "000000000011001001",  -- (p-0.5)^2*pi^2(0.30)=3.917059e-01
    "000000000011000111",  -- (p-0.5)^2*pi^2(0.30)=3.878751e-01
    "000000000011000101",  -- (p-0.5)^2*pi^2(0.30)=3.840631e-01
    "000000000011000011",  -- (p-0.5)^2*pi^2(0.30)=3.802699e-01
    "000000000011000001",  -- (p-0.5)^2*pi^2(0.30)=3.764955e-01
    "000000000010111111",  -- (p-0.5)^2*pi^2(0.31)=3.727400e-01
    "000000000010111101",  -- (p-0.5)^2*pi^2(0.31)=3.690033e-01
    "000000000010111011",  -- (p-0.5)^2*pi^2(0.31)=3.652854e-01
    "000000000010111001",  -- (p-0.5)^2*pi^2(0.31)=3.615863e-01
    "000000000010110111",  -- (p-0.5)^2*pi^2(0.31)=3.579061e-01
    "000000000010110101",  -- (p-0.5)^2*pi^2(0.31)=3.542446e-01
    "000000000010110100",  -- (p-0.5)^2*pi^2(0.31)=3.506020e-01
    "000000000010110010",  -- (p-0.5)^2*pi^2(0.31)=3.469783e-01
    "000000000010110000",  -- (p-0.5)^2*pi^2(0.31)=3.433733e-01
    "000000000010101110",  -- (p-0.5)^2*pi^2(0.31)=3.397872e-01
    "000000000010101100",  -- (p-0.5)^2*pi^2(0.32)=3.362199e-01
    "000000000010101010",  -- (p-0.5)^2*pi^2(0.32)=3.326714e-01
    "000000000010101001",  -- (p-0.5)^2*pi^2(0.32)=3.291418e-01
    "000000000010100111",  -- (p-0.5)^2*pi^2(0.32)=3.256310e-01
    "000000000010100101",  -- (p-0.5)^2*pi^2(0.32)=3.221390e-01
    "000000000010100011",  -- (p-0.5)^2*pi^2(0.32)=3.186658e-01
    "000000000010100001",  -- (p-0.5)^2*pi^2(0.32)=3.152115e-01
    "000000000010100000",  -- (p-0.5)^2*pi^2(0.32)=3.117759e-01
    "000000000010011110",  -- (p-0.5)^2*pi^2(0.32)=3.083593e-01
    "000000000010011100",  -- (p-0.5)^2*pi^2(0.32)=3.049614e-01
    "000000000010011010",  -- (p-0.5)^2*pi^2(0.33)=3.015823e-01
    "000000000010011001",  -- (p-0.5)^2*pi^2(0.33)=2.982221e-01
    "000000000010010111",  -- (p-0.5)^2*pi^2(0.33)=2.948807e-01
    "000000000010010101",  -- (p-0.5)^2*pi^2(0.33)=2.915581e-01
    "000000000010010100",  -- (p-0.5)^2*pi^2(0.33)=2.882544e-01
    "000000000010010010",  -- (p-0.5)^2*pi^2(0.33)=2.849695e-01
    "000000000010010000",  -- (p-0.5)^2*pi^2(0.33)=2.817034e-01
    "000000000010001111",  -- (p-0.5)^2*pi^2(0.33)=2.784561e-01
    "000000000010001101",  -- (p-0.5)^2*pi^2(0.33)=2.752276e-01
    "000000000010001011",  -- (p-0.5)^2*pi^2(0.33)=2.720180e-01
    "000000000010001010",  -- (p-0.5)^2*pi^2(0.33)=2.688272e-01
    "000000000010001000",  -- (p-0.5)^2*pi^2(0.34)=2.656552e-01
    "000000000010000110",  -- (p-0.5)^2*pi^2(0.34)=2.625021e-01
    "000000000010000101",  -- (p-0.5)^2*pi^2(0.34)=2.593678e-01
    "000000000010000011",  -- (p-0.5)^2*pi^2(0.34)=2.562523e-01
    "000000000010000010",  -- (p-0.5)^2*pi^2(0.34)=2.531556e-01
    "000000000010000000",  -- (p-0.5)^2*pi^2(0.34)=2.500777e-01
    "000000000001111110",  -- (p-0.5)^2*pi^2(0.34)=2.470187e-01
    "000000000001111101",  -- (p-0.5)^2*pi^2(0.34)=2.439785e-01
    "000000000001111011",  -- (p-0.5)^2*pi^2(0.34)=2.409571e-01
    "000000000001111010",  -- (p-0.5)^2*pi^2(0.34)=2.379546e-01
    "000000000001111000",  -- (p-0.5)^2*pi^2(0.35)=2.349709e-01
    "000000000001110111",  -- (p-0.5)^2*pi^2(0.35)=2.320060e-01
    "000000000001110101",  -- (p-0.5)^2*pi^2(0.35)=2.290599e-01
    "000000000001110100",  -- (p-0.5)^2*pi^2(0.35)=2.261326e-01
    "000000000001110010",  -- (p-0.5)^2*pi^2(0.35)=2.232242e-01
    "000000000001110001",  -- (p-0.5)^2*pi^2(0.35)=2.203346e-01
    "000000000001101111",  -- (p-0.5)^2*pi^2(0.35)=2.174638e-01
    "000000000001101110",  -- (p-0.5)^2*pi^2(0.35)=2.146119e-01
    "000000000001101100",  -- (p-0.5)^2*pi^2(0.35)=2.117787e-01
    "000000000001101011",  -- (p-0.5)^2*pi^2(0.35)=2.089644e-01
    "000000000001101010",  -- (p-0.5)^2*pi^2(0.36)=2.061690e-01
    "000000000001101000",  -- (p-0.5)^2*pi^2(0.36)=2.033923e-01
    "000000000001100111",  -- (p-0.5)^2*pi^2(0.36)=2.006345e-01
    "000000000001100101",  -- (p-0.5)^2*pi^2(0.36)=1.978955e-01
    "000000000001100100",  -- (p-0.5)^2*pi^2(0.36)=1.951753e-01
    "000000000001100011",  -- (p-0.5)^2*pi^2(0.36)=1.924739e-01
    "000000000001100001",  -- (p-0.5)^2*pi^2(0.36)=1.897914e-01
    "000000000001100000",  -- (p-0.5)^2*pi^2(0.36)=1.871277e-01
    "000000000001011110",  -- (p-0.5)^2*pi^2(0.36)=1.844828e-01
    "000000000001011101",  -- (p-0.5)^2*pi^2(0.36)=1.818568e-01
    "000000000001011100",  -- (p-0.5)^2*pi^2(0.37)=1.792495e-01
    "000000000001011010",  -- (p-0.5)^2*pi^2(0.37)=1.766611e-01
    "000000000001011001",  -- (p-0.5)^2*pi^2(0.37)=1.740915e-01
    "000000000001011000",  -- (p-0.5)^2*pi^2(0.37)=1.715408e-01
    "000000000001010111",  -- (p-0.5)^2*pi^2(0.37)=1.690088e-01
    "000000000001010101",  -- (p-0.5)^2*pi^2(0.37)=1.664957e-01
    "000000000001010100",  -- (p-0.5)^2*pi^2(0.37)=1.640015e-01
    "000000000001010011",  -- (p-0.5)^2*pi^2(0.37)=1.615260e-01
    "000000000001010001",  -- (p-0.5)^2*pi^2(0.37)=1.590694e-01
    "000000000001010000",  -- (p-0.5)^2*pi^2(0.37)=1.566316e-01
    "000000000001001111",  -- (p-0.5)^2*pi^2(0.38)=1.542126e-01
    "000000000001001110",  -- (p-0.5)^2*pi^2(0.38)=1.518124e-01
    "000000000001001101",  -- (p-0.5)^2*pi^2(0.38)=1.494311e-01
    "000000000001001011",  -- (p-0.5)^2*pi^2(0.38)=1.470686e-01
    "000000000001001010",  -- (p-0.5)^2*pi^2(0.38)=1.447249e-01
    "000000000001001001",  -- (p-0.5)^2*pi^2(0.38)=1.424000e-01
    "000000000001001000",  -- (p-0.5)^2*pi^2(0.38)=1.400940e-01
    "000000000001000111",  -- (p-0.5)^2*pi^2(0.38)=1.378068e-01
    "000000000001000101",  -- (p-0.5)^2*pi^2(0.38)=1.355384e-01
    "000000000001000100",  -- (p-0.5)^2*pi^2(0.38)=1.332888e-01
    "000000000001000011",  -- (p-0.5)^2*pi^2(0.38)=1.310581e-01
    "000000000001000010",  -- (p-0.5)^2*pi^2(0.39)=1.288462e-01
    "000000000001000001",  -- (p-0.5)^2*pi^2(0.39)=1.266531e-01
    "000000000001000000",  -- (p-0.5)^2*pi^2(0.39)=1.244788e-01
    "000000000000111111",  -- (p-0.5)^2*pi^2(0.39)=1.223234e-01
    "000000000000111110",  -- (p-0.5)^2*pi^2(0.39)=1.201868e-01
    "000000000000111100",  -- (p-0.5)^2*pi^2(0.39)=1.180690e-01
    "000000000000111011",  -- (p-0.5)^2*pi^2(0.39)=1.159700e-01
    "000000000000111010",  -- (p-0.5)^2*pi^2(0.39)=1.138899e-01
    "000000000000111001",  -- (p-0.5)^2*pi^2(0.39)=1.118286e-01
    "000000000000111000",  -- (p-0.5)^2*pi^2(0.39)=1.097861e-01
    "000000000000110111",  -- (p-0.5)^2*pi^2(0.40)=1.077624e-01
    "000000000000110110",  -- (p-0.5)^2*pi^2(0.40)=1.057576e-01
    "000000000000110101",  -- (p-0.5)^2*pi^2(0.40)=1.037716e-01
    "000000000000110100",  -- (p-0.5)^2*pi^2(0.40)=1.018044e-01
    "000000000000110011",  -- (p-0.5)^2*pi^2(0.40)=9.985603e-02
    "000000000000110010",  -- (p-0.5)^2*pi^2(0.40)=9.792649e-02
    "000000000000110001",  -- (p-0.5)^2*pi^2(0.40)=9.601577e-02
    "000000000000110000",  -- (p-0.5)^2*pi^2(0.40)=9.412388e-02
    "000000000000101111",  -- (p-0.5)^2*pi^2(0.40)=9.225082e-02
    "000000000000101110",  -- (p-0.5)^2*pi^2(0.40)=9.039658e-02
    "000000000000101101",  -- (p-0.5)^2*pi^2(0.41)=8.856116e-02
    "000000000000101100",  -- (p-0.5)^2*pi^2(0.41)=8.674457e-02
    "000000000000101011",  -- (p-0.5)^2*pi^2(0.41)=8.494680e-02
    "000000000000101011",  -- (p-0.5)^2*pi^2(0.41)=8.316786e-02
    "000000000000101010",  -- (p-0.5)^2*pi^2(0.41)=8.140775e-02
    "000000000000101001",  -- (p-0.5)^2*pi^2(0.41)=7.966645e-02
    "000000000000101000",  -- (p-0.5)^2*pi^2(0.41)=7.794399e-02
    "000000000000100111",  -- (p-0.5)^2*pi^2(0.41)=7.624034e-02
    "000000000000100110",  -- (p-0.5)^2*pi^2(0.41)=7.455553e-02
    "000000000000100101",  -- (p-0.5)^2*pi^2(0.41)=7.288953e-02
    "000000000000100100",  -- (p-0.5)^2*pi^2(0.42)=7.124237e-02
    "000000000000100100",  -- (p-0.5)^2*pi^2(0.42)=6.961402e-02
    "000000000000100011",  -- (p-0.5)^2*pi^2(0.42)=6.800450e-02
    "000000000000100010",  -- (p-0.5)^2*pi^2(0.42)=6.641381e-02
    "000000000000100001",  -- (p-0.5)^2*pi^2(0.42)=6.484194e-02
    "000000000000100000",  -- (p-0.5)^2*pi^2(0.42)=6.328890e-02
    "000000000000100000",  -- (p-0.5)^2*pi^2(0.42)=6.175468e-02
    "000000000000011111",  -- (p-0.5)^2*pi^2(0.42)=6.023928e-02
    "000000000000011110",  -- (p-0.5)^2*pi^2(0.42)=5.874271e-02
    "000000000000011101",  -- (p-0.5)^2*pi^2(0.42)=5.726497e-02
    "000000000000011101",  -- (p-0.5)^2*pi^2(0.42)=5.580605e-02
    "000000000000011100",  -- (p-0.5)^2*pi^2(0.43)=5.436595e-02
    "000000000000011011",  -- (p-0.5)^2*pi^2(0.43)=5.294468e-02
    "000000000000011010",  -- (p-0.5)^2*pi^2(0.43)=5.154224e-02
    "000000000000011010",  -- (p-0.5)^2*pi^2(0.43)=5.015862e-02
    "000000000000011001",  -- (p-0.5)^2*pi^2(0.43)=4.879382e-02
    "000000000000011000",  -- (p-0.5)^2*pi^2(0.43)=4.744785e-02
    "000000000000011000",  -- (p-0.5)^2*pi^2(0.43)=4.612070e-02
    "000000000000010111",  -- (p-0.5)^2*pi^2(0.43)=4.481238e-02
    "000000000000010110",  -- (p-0.5)^2*pi^2(0.43)=4.352288e-02
    "000000000000010110",  -- (p-0.5)^2*pi^2(0.43)=4.225221e-02
    "000000000000010101",  -- (p-0.5)^2*pi^2(0.44)=4.100036e-02
    "000000000000010100",  -- (p-0.5)^2*pi^2(0.44)=3.976734e-02
    "000000000000010100",  -- (p-0.5)^2*pi^2(0.44)=3.855314e-02
    "000000000000010011",  -- (p-0.5)^2*pi^2(0.44)=3.735777e-02
    "000000000000010011",  -- (p-0.5)^2*pi^2(0.44)=3.618122e-02
    "000000000000010010",  -- (p-0.5)^2*pi^2(0.44)=3.502350e-02
    "000000000000010001",  -- (p-0.5)^2*pi^2(0.44)=3.388460e-02
    "000000000000010001",  -- (p-0.5)^2*pi^2(0.44)=3.276452e-02
    "000000000000010000",  -- (p-0.5)^2*pi^2(0.44)=3.166327e-02
    "000000000000010000",  -- (p-0.5)^2*pi^2(0.44)=3.058085e-02
    "000000000000001111",  -- (p-0.5)^2*pi^2(0.45)=2.951725e-02
    "000000000000001111",  -- (p-0.5)^2*pi^2(0.45)=2.847247e-02
    "000000000000001110",  -- (p-0.5)^2*pi^2(0.45)=2.744652e-02
    "000000000000001110",  -- (p-0.5)^2*pi^2(0.45)=2.643940e-02
    "000000000000001101",  -- (p-0.5)^2*pi^2(0.45)=2.545110e-02
    "000000000000001101",  -- (p-0.5)^2*pi^2(0.45)=2.448162e-02
    "000000000000001100",  -- (p-0.5)^2*pi^2(0.45)=2.353097e-02
    "000000000000001100",  -- (p-0.5)^2*pi^2(0.45)=2.259914e-02
    "000000000000001011",  -- (p-0.5)^2*pi^2(0.45)=2.168614e-02
    "000000000000001011",  -- (p-0.5)^2*pi^2(0.45)=2.079197e-02
    "000000000000001010",  -- (p-0.5)^2*pi^2(0.46)=1.991661e-02
    "000000000000001010",  -- (p-0.5)^2*pi^2(0.46)=1.906009e-02
    "000000000000001001",  -- (p-0.5)^2*pi^2(0.46)=1.822238e-02
    "000000000000001001",  -- (p-0.5)^2*pi^2(0.46)=1.740351e-02
    "000000000000001001",  -- (p-0.5)^2*pi^2(0.46)=1.660345e-02
    "000000000000001000",  -- (p-0.5)^2*pi^2(0.46)=1.582222e-02
    "000000000000001000",  -- (p-0.5)^2*pi^2(0.46)=1.505982e-02
    "000000000000000111",  -- (p-0.5)^2*pi^2(0.46)=1.431624e-02
    "000000000000000111",  -- (p-0.5)^2*pi^2(0.46)=1.359149e-02
    "000000000000000111",  -- (p-0.5)^2*pi^2(0.46)=1.288556e-02
    "000000000000000110",  -- (p-0.5)^2*pi^2(0.46)=1.219846e-02
    "000000000000000110",  -- (p-0.5)^2*pi^2(0.47)=1.153018e-02
    "000000000000000110",  -- (p-0.5)^2*pi^2(0.47)=1.088072e-02
    "000000000000000101",  -- (p-0.5)^2*pi^2(0.47)=1.025009e-02
    "000000000000000101",  -- (p-0.5)^2*pi^2(0.47)=9.638286e-03
    "000000000000000101",  -- (p-0.5)^2*pi^2(0.47)=9.045305e-03
    "000000000000000100",  -- (p-0.5)^2*pi^2(0.47)=8.471149e-03
    "000000000000000100",  -- (p-0.5)^2*pi^2(0.47)=7.915819e-03
    "000000000000000100",  -- (p-0.5)^2*pi^2(0.47)=7.379312e-03
    "000000000000000100",  -- (p-0.5)^2*pi^2(0.47)=6.861631e-03
    "000000000000000011",  -- (p-0.5)^2*pi^2(0.47)=6.362774e-03
    "000000000000000011",  -- (p-0.5)^2*pi^2(0.48)=5.882743e-03
    "000000000000000011",  -- (p-0.5)^2*pi^2(0.48)=5.421536e-03
    "000000000000000011",  -- (p-0.5)^2*pi^2(0.48)=4.979153e-03
    "000000000000000010",  -- (p-0.5)^2*pi^2(0.48)=4.555596e-03
    "000000000000000010",  -- (p-0.5)^2*pi^2(0.48)=4.150863e-03
    "000000000000000010",  -- (p-0.5)^2*pi^2(0.48)=3.764955e-03
    "000000000000000010",  -- (p-0.5)^2*pi^2(0.48)=3.397872e-03
    "000000000000000010",  -- (p-0.5)^2*pi^2(0.48)=3.049614e-03
    "000000000000000001",  -- (p-0.5)^2*pi^2(0.48)=2.720180e-03
    "000000000000000001",  -- (p-0.5)^2*pi^2(0.48)=2.409571e-03
    "000000000000000001",  -- (p-0.5)^2*pi^2(0.49)=2.117787e-03
    "000000000000000001",  -- (p-0.5)^2*pi^2(0.49)=1.844828e-03
    "000000000000000001",  -- (p-0.5)^2*pi^2(0.49)=1.590694e-03
    "000000000000000001",  -- (p-0.5)^2*pi^2(0.49)=1.355384e-03
    "000000000000000001",  -- (p-0.5)^2*pi^2(0.49)=1.138899e-03
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.49)=9.412388e-04
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.49)=7.624034e-04
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.49)=6.023928e-04
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.49)=4.612070e-04
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.49)=3.388460e-04
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.50)=2.353097e-04
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.50)=1.505982e-04
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.50)=8.471149e-05
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.50)=3.764955e-05
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.50)=9.412388e-06
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.50)=0
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.50)=9.412388e-06
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.50)=3.764955e-05
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.50)=8.471149e-05
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.50)=1.505982e-04
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.50)=2.353097e-04
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.51)=3.388460e-04
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.51)=4.612070e-04
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.51)=6.023928e-04
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.51)=7.624034e-04
    "000000000000000000",  -- (p-0.5)^2*pi^2(0.51)=9.412388e-04
    "000000000000000001",  -- (p-0.5)^2*pi^2(0.51)=1.138899e-03
    "000000000000000001",  -- (p-0.5)^2*pi^2(0.51)=1.355384e-03
    "000000000000000001",  -- (p-0.5)^2*pi^2(0.51)=1.590694e-03
    "000000000000000001",  -- (p-0.5)^2*pi^2(0.51)=1.844828e-03
    "000000000000000001",  -- (p-0.5)^2*pi^2(0.51)=2.117787e-03
    "000000000000000001",  -- (p-0.5)^2*pi^2(0.52)=2.409571e-03
    "000000000000000001",  -- (p-0.5)^2*pi^2(0.52)=2.720180e-03
    "000000000000000010",  -- (p-0.5)^2*pi^2(0.52)=3.049614e-03
    "000000000000000010",  -- (p-0.5)^2*pi^2(0.52)=3.397872e-03
    "000000000000000010",  -- (p-0.5)^2*pi^2(0.52)=3.764955e-03
    "000000000000000010",  -- (p-0.5)^2*pi^2(0.52)=4.150863e-03
    "000000000000000010",  -- (p-0.5)^2*pi^2(0.52)=4.555596e-03
    "000000000000000011",  -- (p-0.5)^2*pi^2(0.52)=4.979153e-03
    "000000000000000011",  -- (p-0.5)^2*pi^2(0.52)=5.421536e-03
    "000000000000000011",  -- (p-0.5)^2*pi^2(0.52)=5.882743e-03
    "000000000000000011",  -- (p-0.5)^2*pi^2(0.53)=6.362774e-03
    "000000000000000100",  -- (p-0.5)^2*pi^2(0.53)=6.861631e-03
    "000000000000000100",  -- (p-0.5)^2*pi^2(0.53)=7.379312e-03
    "000000000000000100",  -- (p-0.5)^2*pi^2(0.53)=7.915819e-03
    "000000000000000100",  -- (p-0.5)^2*pi^2(0.53)=8.471149e-03
    "000000000000000101",  -- (p-0.5)^2*pi^2(0.53)=9.045305e-03
    "000000000000000101",  -- (p-0.5)^2*pi^2(0.53)=9.638286e-03
    "000000000000000101",  -- (p-0.5)^2*pi^2(0.53)=1.025009e-02
    "000000000000000110",  -- (p-0.5)^2*pi^2(0.53)=1.088072e-02
    "000000000000000110",  -- (p-0.5)^2*pi^2(0.53)=1.153018e-02
    "000000000000000110",  -- (p-0.5)^2*pi^2(0.54)=1.219846e-02
    "000000000000000111",  -- (p-0.5)^2*pi^2(0.54)=1.288556e-02
    "000000000000000111",  -- (p-0.5)^2*pi^2(0.54)=1.359149e-02
    "000000000000000111",  -- (p-0.5)^2*pi^2(0.54)=1.431624e-02
    "000000000000001000",  -- (p-0.5)^2*pi^2(0.54)=1.505982e-02
    "000000000000001000",  -- (p-0.5)^2*pi^2(0.54)=1.582222e-02
    "000000000000001001",  -- (p-0.5)^2*pi^2(0.54)=1.660345e-02
    "000000000000001001",  -- (p-0.5)^2*pi^2(0.54)=1.740351e-02
    "000000000000001001",  -- (p-0.5)^2*pi^2(0.54)=1.822238e-02
    "000000000000001010",  -- (p-0.5)^2*pi^2(0.54)=1.906009e-02
    "000000000000001010",  -- (p-0.5)^2*pi^2(0.54)=1.991661e-02
    "000000000000001011",  -- (p-0.5)^2*pi^2(0.55)=2.079197e-02
    "000000000000001011",  -- (p-0.5)^2*pi^2(0.55)=2.168614e-02
    "000000000000001100",  -- (p-0.5)^2*pi^2(0.55)=2.259914e-02
    "000000000000001100",  -- (p-0.5)^2*pi^2(0.55)=2.353097e-02
    "000000000000001101",  -- (p-0.5)^2*pi^2(0.55)=2.448162e-02
    "000000000000001101",  -- (p-0.5)^2*pi^2(0.55)=2.545110e-02
    "000000000000001110",  -- (p-0.5)^2*pi^2(0.55)=2.643940e-02
    "000000000000001110",  -- (p-0.5)^2*pi^2(0.55)=2.744652e-02
    "000000000000001111",  -- (p-0.5)^2*pi^2(0.55)=2.847247e-02
    "000000000000001111",  -- (p-0.5)^2*pi^2(0.55)=2.951725e-02
    "000000000000010000",  -- (p-0.5)^2*pi^2(0.56)=3.058085e-02
    "000000000000010000",  -- (p-0.5)^2*pi^2(0.56)=3.166327e-02
    "000000000000010001",  -- (p-0.5)^2*pi^2(0.56)=3.276452e-02
    "000000000000010001",  -- (p-0.5)^2*pi^2(0.56)=3.388460e-02
    "000000000000010010",  -- (p-0.5)^2*pi^2(0.56)=3.502350e-02
    "000000000000010011",  -- (p-0.5)^2*pi^2(0.56)=3.618122e-02
    "000000000000010011",  -- (p-0.5)^2*pi^2(0.56)=3.735777e-02
    "000000000000010100",  -- (p-0.5)^2*pi^2(0.56)=3.855314e-02
    "000000000000010100",  -- (p-0.5)^2*pi^2(0.56)=3.976734e-02
    "000000000000010101",  -- (p-0.5)^2*pi^2(0.56)=4.100036e-02
    "000000000000010110",  -- (p-0.5)^2*pi^2(0.57)=4.225221e-02
    "000000000000010110",  -- (p-0.5)^2*pi^2(0.57)=4.352288e-02
    "000000000000010111",  -- (p-0.5)^2*pi^2(0.57)=4.481238e-02
    "000000000000011000",  -- (p-0.5)^2*pi^2(0.57)=4.612070e-02
    "000000000000011000",  -- (p-0.5)^2*pi^2(0.57)=4.744785e-02
    "000000000000011001",  -- (p-0.5)^2*pi^2(0.57)=4.879382e-02
    "000000000000011010",  -- (p-0.5)^2*pi^2(0.57)=5.015862e-02
    "000000000000011010",  -- (p-0.5)^2*pi^2(0.57)=5.154224e-02
    "000000000000011011",  -- (p-0.5)^2*pi^2(0.57)=5.294468e-02
    "000000000000011100",  -- (p-0.5)^2*pi^2(0.57)=5.436595e-02
    "000000000000011101",  -- (p-0.5)^2*pi^2(0.58)=5.580605e-02
    "000000000000011101",  -- (p-0.5)^2*pi^2(0.58)=5.726497e-02
    "000000000000011110",  -- (p-0.5)^2*pi^2(0.58)=5.874271e-02
    "000000000000011111",  -- (p-0.5)^2*pi^2(0.58)=6.023928e-02
    "000000000000100000",  -- (p-0.5)^2*pi^2(0.58)=6.175468e-02
    "000000000000100000",  -- (p-0.5)^2*pi^2(0.58)=6.328890e-02
    "000000000000100001",  -- (p-0.5)^2*pi^2(0.58)=6.484194e-02
    "000000000000100010",  -- (p-0.5)^2*pi^2(0.58)=6.641381e-02
    "000000000000100011",  -- (p-0.5)^2*pi^2(0.58)=6.800450e-02
    "000000000000100100",  -- (p-0.5)^2*pi^2(0.58)=6.961402e-02
    "000000000000100100",  -- (p-0.5)^2*pi^2(0.58)=7.124237e-02
    "000000000000100101",  -- (p-0.5)^2*pi^2(0.59)=7.288953e-02
    "000000000000100110",  -- (p-0.5)^2*pi^2(0.59)=7.455553e-02
    "000000000000100111",  -- (p-0.5)^2*pi^2(0.59)=7.624034e-02
    "000000000000101000",  -- (p-0.5)^2*pi^2(0.59)=7.794399e-02
    "000000000000101001",  -- (p-0.5)^2*pi^2(0.59)=7.966645e-02
    "000000000000101010",  -- (p-0.5)^2*pi^2(0.59)=8.140775e-02
    "000000000000101011",  -- (p-0.5)^2*pi^2(0.59)=8.316786e-02
    "000000000000101011",  -- (p-0.5)^2*pi^2(0.59)=8.494680e-02
    "000000000000101100",  -- (p-0.5)^2*pi^2(0.59)=8.674457e-02
    "000000000000101101",  -- (p-0.5)^2*pi^2(0.59)=8.856116e-02
    "000000000000101110",  -- (p-0.5)^2*pi^2(0.60)=9.039658e-02
    "000000000000101111",  -- (p-0.5)^2*pi^2(0.60)=9.225082e-02
    "000000000000110000",  -- (p-0.5)^2*pi^2(0.60)=9.412388e-02
    "000000000000110001",  -- (p-0.5)^2*pi^2(0.60)=9.601577e-02
    "000000000000110010",  -- (p-0.5)^2*pi^2(0.60)=9.792649e-02
    "000000000000110011",  -- (p-0.5)^2*pi^2(0.60)=9.985603e-02
    "000000000000110100",  -- (p-0.5)^2*pi^2(0.60)=1.018044e-01
    "000000000000110101",  -- (p-0.5)^2*pi^2(0.60)=1.037716e-01
    "000000000000110110",  -- (p-0.5)^2*pi^2(0.60)=1.057576e-01
    "000000000000110111",  -- (p-0.5)^2*pi^2(0.60)=1.077624e-01
    "000000000000111000",  -- (p-0.5)^2*pi^2(0.61)=1.097861e-01
    "000000000000111001",  -- (p-0.5)^2*pi^2(0.61)=1.118286e-01
    "000000000000111010",  -- (p-0.5)^2*pi^2(0.61)=1.138899e-01
    "000000000000111011",  -- (p-0.5)^2*pi^2(0.61)=1.159700e-01
    "000000000000111100",  -- (p-0.5)^2*pi^2(0.61)=1.180690e-01
    "000000000000111110",  -- (p-0.5)^2*pi^2(0.61)=1.201868e-01
    "000000000000111111",  -- (p-0.5)^2*pi^2(0.61)=1.223234e-01
    "000000000001000000",  -- (p-0.5)^2*pi^2(0.61)=1.244788e-01
    "000000000001000001",  -- (p-0.5)^2*pi^2(0.61)=1.266531e-01
    "000000000001000010",  -- (p-0.5)^2*pi^2(0.61)=1.288462e-01
    "000000000001000011",  -- (p-0.5)^2*pi^2(0.62)=1.310581e-01
    "000000000001000100",  -- (p-0.5)^2*pi^2(0.62)=1.332888e-01
    "000000000001000101",  -- (p-0.5)^2*pi^2(0.62)=1.355384e-01
    "000000000001000111",  -- (p-0.5)^2*pi^2(0.62)=1.378068e-01
    "000000000001001000",  -- (p-0.5)^2*pi^2(0.62)=1.400940e-01
    "000000000001001001",  -- (p-0.5)^2*pi^2(0.62)=1.424000e-01
    "000000000001001010",  -- (p-0.5)^2*pi^2(0.62)=1.447249e-01
    "000000000001001011",  -- (p-0.5)^2*pi^2(0.62)=1.470686e-01
    "000000000001001101",  -- (p-0.5)^2*pi^2(0.62)=1.494311e-01
    "000000000001001110",  -- (p-0.5)^2*pi^2(0.62)=1.518124e-01
    "000000000001001111",  -- (p-0.5)^2*pi^2(0.62)=1.542126e-01
    "000000000001010000",  -- (p-0.5)^2*pi^2(0.63)=1.566316e-01
    "000000000001010001",  -- (p-0.5)^2*pi^2(0.63)=1.590694e-01
    "000000000001010011",  -- (p-0.5)^2*pi^2(0.63)=1.615260e-01
    "000000000001010100",  -- (p-0.5)^2*pi^2(0.63)=1.640015e-01
    "000000000001010101",  -- (p-0.5)^2*pi^2(0.63)=1.664957e-01
    "000000000001010111",  -- (p-0.5)^2*pi^2(0.63)=1.690088e-01
    "000000000001011000",  -- (p-0.5)^2*pi^2(0.63)=1.715408e-01
    "000000000001011001",  -- (p-0.5)^2*pi^2(0.63)=1.740915e-01
    "000000000001011010",  -- (p-0.5)^2*pi^2(0.63)=1.766611e-01
    "000000000001011100",  -- (p-0.5)^2*pi^2(0.63)=1.792495e-01
    "000000000001011101",  -- (p-0.5)^2*pi^2(0.64)=1.818568e-01
    "000000000001011110",  -- (p-0.5)^2*pi^2(0.64)=1.844828e-01
    "000000000001100000",  -- (p-0.5)^2*pi^2(0.64)=1.871277e-01
    "000000000001100001",  -- (p-0.5)^2*pi^2(0.64)=1.897914e-01
    "000000000001100011",  -- (p-0.5)^2*pi^2(0.64)=1.924739e-01
    "000000000001100100",  -- (p-0.5)^2*pi^2(0.64)=1.951753e-01
    "000000000001100101",  -- (p-0.5)^2*pi^2(0.64)=1.978955e-01
    "000000000001100111",  -- (p-0.5)^2*pi^2(0.64)=2.006345e-01
    "000000000001101000",  -- (p-0.5)^2*pi^2(0.64)=2.033923e-01
    "000000000001101010",  -- (p-0.5)^2*pi^2(0.64)=2.061690e-01
    "000000000001101011",  -- (p-0.5)^2*pi^2(0.65)=2.089644e-01
    "000000000001101100",  -- (p-0.5)^2*pi^2(0.65)=2.117787e-01
    "000000000001101110",  -- (p-0.5)^2*pi^2(0.65)=2.146119e-01
    "000000000001101111",  -- (p-0.5)^2*pi^2(0.65)=2.174638e-01
    "000000000001110001",  -- (p-0.5)^2*pi^2(0.65)=2.203346e-01
    "000000000001110010",  -- (p-0.5)^2*pi^2(0.65)=2.232242e-01
    "000000000001110100",  -- (p-0.5)^2*pi^2(0.65)=2.261326e-01
    "000000000001110101",  -- (p-0.5)^2*pi^2(0.65)=2.290599e-01
    "000000000001110111",  -- (p-0.5)^2*pi^2(0.65)=2.320060e-01
    "000000000001111000",  -- (p-0.5)^2*pi^2(0.65)=2.349709e-01
    "000000000001111010",  -- (p-0.5)^2*pi^2(0.66)=2.379546e-01
    "000000000001111011",  -- (p-0.5)^2*pi^2(0.66)=2.409571e-01
    "000000000001111101",  -- (p-0.5)^2*pi^2(0.66)=2.439785e-01
    "000000000001111110",  -- (p-0.5)^2*pi^2(0.66)=2.470187e-01
    "000000000010000000",  -- (p-0.5)^2*pi^2(0.66)=2.500777e-01
    "000000000010000010",  -- (p-0.5)^2*pi^2(0.66)=2.531556e-01
    "000000000010000011",  -- (p-0.5)^2*pi^2(0.66)=2.562523e-01
    "000000000010000101",  -- (p-0.5)^2*pi^2(0.66)=2.593678e-01
    "000000000010000110",  -- (p-0.5)^2*pi^2(0.66)=2.625021e-01
    "000000000010001000",  -- (p-0.5)^2*pi^2(0.66)=2.656552e-01
    "000000000010001010",  -- (p-0.5)^2*pi^2(0.67)=2.688272e-01
    "000000000010001011",  -- (p-0.5)^2*pi^2(0.67)=2.720180e-01
    "000000000010001101",  -- (p-0.5)^2*pi^2(0.67)=2.752276e-01
    "000000000010001111",  -- (p-0.5)^2*pi^2(0.67)=2.784561e-01
    "000000000010010000",  -- (p-0.5)^2*pi^2(0.67)=2.817034e-01
    "000000000010010010",  -- (p-0.5)^2*pi^2(0.67)=2.849695e-01
    "000000000010010100",  -- (p-0.5)^2*pi^2(0.67)=2.882544e-01
    "000000000010010101",  -- (p-0.5)^2*pi^2(0.67)=2.915581e-01
    "000000000010010111",  -- (p-0.5)^2*pi^2(0.67)=2.948807e-01
    "000000000010011001",  -- (p-0.5)^2*pi^2(0.67)=2.982221e-01
    "000000000010011010",  -- (p-0.5)^2*pi^2(0.67)=3.015823e-01
    "000000000010011100",  -- (p-0.5)^2*pi^2(0.68)=3.049614e-01
    "000000000010011110",  -- (p-0.5)^2*pi^2(0.68)=3.083593e-01
    "000000000010100000",  -- (p-0.5)^2*pi^2(0.68)=3.117759e-01
    "000000000010100001",  -- (p-0.5)^2*pi^2(0.68)=3.152115e-01
    "000000000010100011",  -- (p-0.5)^2*pi^2(0.68)=3.186658e-01
    "000000000010100101",  -- (p-0.5)^2*pi^2(0.68)=3.221390e-01
    "000000000010100111",  -- (p-0.5)^2*pi^2(0.68)=3.256310e-01
    "000000000010101001",  -- (p-0.5)^2*pi^2(0.68)=3.291418e-01
    "000000000010101010",  -- (p-0.5)^2*pi^2(0.68)=3.326714e-01
    "000000000010101100",  -- (p-0.5)^2*pi^2(0.68)=3.362199e-01
    "000000000010101110",  -- (p-0.5)^2*pi^2(0.69)=3.397872e-01
    "000000000010110000",  -- (p-0.5)^2*pi^2(0.69)=3.433733e-01
    "000000000010110010",  -- (p-0.5)^2*pi^2(0.69)=3.469783e-01
    "000000000010110100",  -- (p-0.5)^2*pi^2(0.69)=3.506020e-01
    "000000000010110101",  -- (p-0.5)^2*pi^2(0.69)=3.542446e-01
    "000000000010110111",  -- (p-0.5)^2*pi^2(0.69)=3.579061e-01
    "000000000010111001",  -- (p-0.5)^2*pi^2(0.69)=3.615863e-01
    "000000000010111011",  -- (p-0.5)^2*pi^2(0.69)=3.652854e-01
    "000000000010111101",  -- (p-0.5)^2*pi^2(0.69)=3.690033e-01
    "000000000010111111",  -- (p-0.5)^2*pi^2(0.69)=3.727400e-01
    "000000000011000001",  -- (p-0.5)^2*pi^2(0.70)=3.764955e-01
    "000000000011000011",  -- (p-0.5)^2*pi^2(0.70)=3.802699e-01
    "000000000011000101",  -- (p-0.5)^2*pi^2(0.70)=3.840631e-01
    "000000000011000111",  -- (p-0.5)^2*pi^2(0.70)=3.878751e-01
    "000000000011001001",  -- (p-0.5)^2*pi^2(0.70)=3.917059e-01
    "000000000011001011",  -- (p-0.5)^2*pi^2(0.70)=3.955556e-01
    "000000000011001101",  -- (p-0.5)^2*pi^2(0.70)=3.994241e-01
    "000000000011001110",  -- (p-0.5)^2*pi^2(0.70)=4.033114e-01
    "000000000011010000",  -- (p-0.5)^2*pi^2(0.70)=4.072176e-01
    "000000000011010011",  -- (p-0.5)^2*pi^2(0.70)=4.111425e-01
    "000000000011010101",  -- (p-0.5)^2*pi^2(0.71)=4.150863e-01
    "000000000011010111",  -- (p-0.5)^2*pi^2(0.71)=4.190489e-01
    "000000000011011001",  -- (p-0.5)^2*pi^2(0.71)=4.230304e-01
    "000000000011011011",  -- (p-0.5)^2*pi^2(0.71)=4.270306e-01
    "000000000011011101",  -- (p-0.5)^2*pi^2(0.71)=4.310497e-01
    "000000000011011111",  -- (p-0.5)^2*pi^2(0.71)=4.350876e-01
    "000000000011100001",  -- (p-0.5)^2*pi^2(0.71)=4.391444e-01
    "000000000011100011",  -- (p-0.5)^2*pi^2(0.71)=4.432199e-01
    "000000000011100101",  -- (p-0.5)^2*pi^2(0.71)=4.473143e-01
    "000000000011100111",  -- (p-0.5)^2*pi^2(0.71)=4.514276e-01
    "000000000011101001",  -- (p-0.5)^2*pi^2(0.71)=4.555596e-01
    "000000000011101011",  -- (p-0.5)^2*pi^2(0.72)=4.597105e-01
    "000000000011101110",  -- (p-0.5)^2*pi^2(0.72)=4.638801e-01
    "000000000011110000",  -- (p-0.5)^2*pi^2(0.72)=4.680687e-01
    "000000000011110010",  -- (p-0.5)^2*pi^2(0.72)=4.722760e-01
    "000000000011110100",  -- (p-0.5)^2*pi^2(0.72)=4.765022e-01
    "000000000011110110",  -- (p-0.5)^2*pi^2(0.72)=4.807471e-01
    "000000000011111000",  -- (p-0.5)^2*pi^2(0.72)=4.850110e-01
    "000000000011111011",  -- (p-0.5)^2*pi^2(0.72)=4.892936e-01
    "000000000011111101",  -- (p-0.5)^2*pi^2(0.72)=4.935951e-01
    "000000000011111111",  -- (p-0.5)^2*pi^2(0.72)=4.979153e-01
    "000000000100000001",  -- (p-0.5)^2*pi^2(0.73)=5.022544e-01
    "000000000100000011",  -- (p-0.5)^2*pi^2(0.73)=5.066124e-01
    "000000000100000110",  -- (p-0.5)^2*pi^2(0.73)=5.109891e-01
    "000000000100001000",  -- (p-0.5)^2*pi^2(0.73)=5.153847e-01
    "000000000100001010",  -- (p-0.5)^2*pi^2(0.73)=5.197991e-01
    "000000000100001100",  -- (p-0.5)^2*pi^2(0.73)=5.242324e-01
    "000000000100001111",  -- (p-0.5)^2*pi^2(0.73)=5.286844e-01
    "000000000100010001",  -- (p-0.5)^2*pi^2(0.73)=5.331553e-01
    "000000000100010011",  -- (p-0.5)^2*pi^2(0.73)=5.376450e-01
    "000000000100010110",  -- (p-0.5)^2*pi^2(0.73)=5.421536e-01
    "000000000100011000",  -- (p-0.5)^2*pi^2(0.74)=5.466809e-01
    "000000000100011010",  -- (p-0.5)^2*pi^2(0.74)=5.512271e-01
    "000000000100011101",  -- (p-0.5)^2*pi^2(0.74)=5.557921e-01
    "000000000100011111",  -- (p-0.5)^2*pi^2(0.74)=5.603759e-01
    "000000000100100001",  -- (p-0.5)^2*pi^2(0.74)=5.649786e-01
    "000000000100100100",  -- (p-0.5)^2*pi^2(0.74)=5.696001e-01
    "000000000100100110",  -- (p-0.5)^2*pi^2(0.74)=5.742404e-01
    "000000000100101000",  -- (p-0.5)^2*pi^2(0.74)=5.788995e-01
    "000000000100101011",  -- (p-0.5)^2*pi^2(0.74)=5.835775e-01
    "000000000100101101",  -- (p-0.5)^2*pi^2(0.74)=5.882743e-01
    "000000000100110000",  -- (p-0.5)^2*pi^2(0.75)=5.929899e-01
    "000000000100110010",  -- (p-0.5)^2*pi^2(0.75)=5.977243e-01
    "000000000100110100",  -- (p-0.5)^2*pi^2(0.75)=6.024776e-01
    "000000000100110111",  -- (p-0.5)^2*pi^2(0.75)=6.072496e-01
    "000000000100111001",  -- (p-0.5)^2*pi^2(0.75)=6.120405e-01
    "000000000100111100",  -- (p-0.5)^2*pi^2(0.75)=6.168503e-01
    "000000000100111110",  -- (p-0.5)^2*pi^2(0.75)=6.216788e-01
    "000000000101000001",  -- (p-0.5)^2*pi^2(0.75)=6.265262e-01
    "000000000101000011",  -- (p-0.5)^2*pi^2(0.75)=6.313924e-01
    "000000000101000110",  -- (p-0.5)^2*pi^2(0.75)=6.362774e-01
    "000000000101001000",  -- (p-0.5)^2*pi^2(0.75)=6.411813e-01
    "000000000101001011",  -- (p-0.5)^2*pi^2(0.76)=6.461040e-01
    "000000000101001101",  -- (p-0.5)^2*pi^2(0.76)=6.510455e-01
    "000000000101010000",  -- (p-0.5)^2*pi^2(0.76)=6.560058e-01
    "000000000101010010",  -- (p-0.5)^2*pi^2(0.76)=6.609850e-01
    "000000000101010101",  -- (p-0.5)^2*pi^2(0.76)=6.659829e-01
    "000000000101011000",  -- (p-0.5)^2*pi^2(0.76)=6.709997e-01
    "000000000101011010",  -- (p-0.5)^2*pi^2(0.76)=6.760354e-01
    "000000000101011101",  -- (p-0.5)^2*pi^2(0.76)=6.810898e-01
    "000000000101011111",  -- (p-0.5)^2*pi^2(0.76)=6.861631e-01
    "000000000101100010",  -- (p-0.5)^2*pi^2(0.76)=6.912552e-01
    "000000000101100101",  -- (p-0.5)^2*pi^2(0.77)=6.963661e-01
    "000000000101100111",  -- (p-0.5)^2*pi^2(0.77)=7.014959e-01
    "000000000101101010",  -- (p-0.5)^2*pi^2(0.77)=7.066445e-01
    "000000000101101100",  -- (p-0.5)^2*pi^2(0.77)=7.118119e-01
    "000000000101101111",  -- (p-0.5)^2*pi^2(0.77)=7.169981e-01
    "000000000101110010",  -- (p-0.5)^2*pi^2(0.77)=7.222031e-01
    "000000000101110100",  -- (p-0.5)^2*pi^2(0.77)=7.274270e-01
    "000000000101110111",  -- (p-0.5)^2*pi^2(0.77)=7.326697e-01
    "000000000101111010",  -- (p-0.5)^2*pi^2(0.77)=7.379312e-01
    "000000000101111101",  -- (p-0.5)^2*pi^2(0.77)=7.432116e-01
    "000000000101111111",  -- (p-0.5)^2*pi^2(0.78)=7.485108e-01
    "000000000110000010",  -- (p-0.5)^2*pi^2(0.78)=7.538288e-01
    "000000000110000101",  -- (p-0.5)^2*pi^2(0.78)=7.591656e-01
    "000000000110000111",  -- (p-0.5)^2*pi^2(0.78)=7.645212e-01
    "000000000110001010",  -- (p-0.5)^2*pi^2(0.78)=7.698957e-01
    "000000000110001101",  -- (p-0.5)^2*pi^2(0.78)=7.752890e-01
    "000000000110010000",  -- (p-0.5)^2*pi^2(0.78)=7.807011e-01
    "000000000110010010",  -- (p-0.5)^2*pi^2(0.78)=7.861321e-01
    "000000000110010101",  -- (p-0.5)^2*pi^2(0.78)=7.915819e-01
    "000000000110011000",  -- (p-0.5)^2*pi^2(0.78)=7.970504e-01
    "000000000110011011",  -- (p-0.5)^2*pi^2(0.79)=8.025379e-01
    "000000000110011110",  -- (p-0.5)^2*pi^2(0.79)=8.080441e-01
    "000000000110100001",  -- (p-0.5)^2*pi^2(0.79)=8.135692e-01
    "000000000110100011",  -- (p-0.5)^2*pi^2(0.79)=8.191131e-01
    "000000000110100110",  -- (p-0.5)^2*pi^2(0.79)=8.246758e-01
    "000000000110101001",  -- (p-0.5)^2*pi^2(0.79)=8.302574e-01
    "000000000110101100",  -- (p-0.5)^2*pi^2(0.79)=8.358577e-01
    "000000000110101111",  -- (p-0.5)^2*pi^2(0.79)=8.414769e-01
    "000000000110110010",  -- (p-0.5)^2*pi^2(0.79)=8.471149e-01
    "000000000110110101",  -- (p-0.5)^2*pi^2(0.79)=8.527718e-01
    "000000000110111000",  -- (p-0.5)^2*pi^2(0.79)=8.584475e-01
    "000000000110111010",  -- (p-0.5)^2*pi^2(0.80)=8.641420e-01
    "000000000110111101",  -- (p-0.5)^2*pi^2(0.80)=8.698553e-01
    "000000000111000000",  -- (p-0.5)^2*pi^2(0.80)=8.755874e-01
    "000000000111000011",  -- (p-0.5)^2*pi^2(0.80)=8.813384e-01
    "000000000111000110",  -- (p-0.5)^2*pi^2(0.80)=8.871082e-01
    "000000000111001001",  -- (p-0.5)^2*pi^2(0.80)=8.928968e-01
    "000000000111001100",  -- (p-0.5)^2*pi^2(0.80)=8.987042e-01
    "000000000111001111",  -- (p-0.5)^2*pi^2(0.80)=9.045305e-01
    "000000000111010010",  -- (p-0.5)^2*pi^2(0.80)=9.103756e-01
    "000000000111010101",  -- (p-0.5)^2*pi^2(0.80)=9.162395e-01
    "000000000111011000",  -- (p-0.5)^2*pi^2(0.81)=9.221223e-01
    "000000000111011011",  -- (p-0.5)^2*pi^2(0.81)=9.280238e-01
    "000000000111011110",  -- (p-0.5)^2*pi^2(0.81)=9.339442e-01
    "000000000111100001",  -- (p-0.5)^2*pi^2(0.81)=9.398834e-01
    "000000000111100100",  -- (p-0.5)^2*pi^2(0.81)=9.458415e-01
    "000000000111100111",  -- (p-0.5)^2*pi^2(0.81)=9.518183e-01
    "000000000111101010",  -- (p-0.5)^2*pi^2(0.81)=9.578140e-01
    "000000000111101101",  -- (p-0.5)^2*pi^2(0.81)=9.638286e-01
    "000000000111110001",  -- (p-0.5)^2*pi^2(0.81)=9.698619e-01
    "000000000111110100",  -- (p-0.5)^2*pi^2(0.81)=9.759141e-01
    "000000000111110111",  -- (p-0.5)^2*pi^2(0.82)=9.819851e-01
    "000000000111111010",  -- (p-0.5)^2*pi^2(0.82)=9.880749e-01
    "000000000111111101",  -- (p-0.5)^2*pi^2(0.82)=9.941835e-01
    "000000001000000000",  -- (p-0.5)^2*pi^2(0.82)=1.000311e+00
    "000000001000000011",  -- (p-0.5)^2*pi^2(0.82)=1.006457e+00
    "000000001000000110",  -- (p-0.5)^2*pi^2(0.82)=1.012622e+00
    "000000001000001010",  -- (p-0.5)^2*pi^2(0.82)=1.018806e+00
    "000000001000001101",  -- (p-0.5)^2*pi^2(0.82)=1.025009e+00
    "000000001000010000",  -- (p-0.5)^2*pi^2(0.82)=1.031231e+00
    "000000001000010011",  -- (p-0.5)^2*pi^2(0.82)=1.037471e+00
    "000000001000010110",  -- (p-0.5)^2*pi^2(0.83)=1.043730e+00
    "000000001000011010",  -- (p-0.5)^2*pi^2(0.83)=1.050008e+00
    "000000001000011101",  -- (p-0.5)^2*pi^2(0.83)=1.056305e+00
    "000000001000100000",  -- (p-0.5)^2*pi^2(0.83)=1.062621e+00
    "000000001000100011",  -- (p-0.5)^2*pi^2(0.83)=1.068956e+00
    "000000001000100111",  -- (p-0.5)^2*pi^2(0.83)=1.075309e+00
    "000000001000101010",  -- (p-0.5)^2*pi^2(0.83)=1.081681e+00
    "000000001000101101",  -- (p-0.5)^2*pi^2(0.83)=1.088072e+00
    "000000001000110000",  -- (p-0.5)^2*pi^2(0.83)=1.094482e+00
    "000000001000110100",  -- (p-0.5)^2*pi^2(0.83)=1.100911e+00
    "000000001000110111",  -- (p-0.5)^2*pi^2(0.83)=1.107358e+00
    "000000001000111010",  -- (p-0.5)^2*pi^2(0.84)=1.113824e+00
    "000000001000111110",  -- (p-0.5)^2*pi^2(0.84)=1.120310e+00
    "000000001001000001",  -- (p-0.5)^2*pi^2(0.84)=1.126813e+00
    "000000001001000100",  -- (p-0.5)^2*pi^2(0.84)=1.133336e+00
    "000000001001001000",  -- (p-0.5)^2*pi^2(0.84)=1.139878e+00
    "000000001001001011",  -- (p-0.5)^2*pi^2(0.84)=1.146438e+00
    "000000001001001110",  -- (p-0.5)^2*pi^2(0.84)=1.153018e+00
    "000000001001010010",  -- (p-0.5)^2*pi^2(0.84)=1.159616e+00
    "000000001001010101",  -- (p-0.5)^2*pi^2(0.84)=1.166233e+00
    "000000001001011001",  -- (p-0.5)^2*pi^2(0.84)=1.172868e+00
    "000000001001011100",  -- (p-0.5)^2*pi^2(0.85)=1.179523e+00
    "000000001001011111",  -- (p-0.5)^2*pi^2(0.85)=1.186196e+00
    "000000001001100011",  -- (p-0.5)^2*pi^2(0.85)=1.192888e+00
    "000000001001100110",  -- (p-0.5)^2*pi^2(0.85)=1.199599e+00
    "000000001001101010",  -- (p-0.5)^2*pi^2(0.85)=1.206329e+00
    "000000001001101101",  -- (p-0.5)^2*pi^2(0.85)=1.213078e+00
    "000000001001110001",  -- (p-0.5)^2*pi^2(0.85)=1.219846e+00
    "000000001001110100",  -- (p-0.5)^2*pi^2(0.85)=1.226632e+00
    "000000001001111000",  -- (p-0.5)^2*pi^2(0.85)=1.233437e+00
    "000000001001111011",  -- (p-0.5)^2*pi^2(0.85)=1.240261e+00
    "000000001001111111",  -- (p-0.5)^2*pi^2(0.86)=1.247104e+00
    "000000001010000010",  -- (p-0.5)^2*pi^2(0.86)=1.253965e+00
    "000000001010000110",  -- (p-0.5)^2*pi^2(0.86)=1.260846e+00
    "000000001010001001",  -- (p-0.5)^2*pi^2(0.86)=1.267745e+00
    "000000001010001101",  -- (p-0.5)^2*pi^2(0.86)=1.274663e+00
    "000000001010010000",  -- (p-0.5)^2*pi^2(0.86)=1.281600e+00
    "000000001010010100",  -- (p-0.5)^2*pi^2(0.86)=1.288556e+00
    "000000001010010111",  -- (p-0.5)^2*pi^2(0.86)=1.295531e+00
    "000000001010011011",  -- (p-0.5)^2*pi^2(0.86)=1.302524e+00
    "000000001010011110",  -- (p-0.5)^2*pi^2(0.86)=1.309536e+00
    "000000001010100010",  -- (p-0.5)^2*pi^2(0.87)=1.316567e+00
    "000000001010100110",  -- (p-0.5)^2*pi^2(0.87)=1.323617e+00
    "000000001010101001",  -- (p-0.5)^2*pi^2(0.87)=1.330686e+00
    "000000001010101101",  -- (p-0.5)^2*pi^2(0.87)=1.337773e+00
    "000000001010110001",  -- (p-0.5)^2*pi^2(0.87)=1.344880e+00
    "000000001010110100",  -- (p-0.5)^2*pi^2(0.87)=1.352005e+00
    "000000001010111000",  -- (p-0.5)^2*pi^2(0.87)=1.359149e+00
    "000000001010111100",  -- (p-0.5)^2*pi^2(0.87)=1.366312e+00
    "000000001010111111",  -- (p-0.5)^2*pi^2(0.87)=1.373493e+00
    "000000001011000011",  -- (p-0.5)^2*pi^2(0.87)=1.380694e+00
    "000000001011000111",  -- (p-0.5)^2*pi^2(0.88)=1.387913e+00
    "000000001011001010",  -- (p-0.5)^2*pi^2(0.88)=1.395151e+00
    "000000001011001110",  -- (p-0.5)^2*pi^2(0.88)=1.402408e+00
    "000000001011010010",  -- (p-0.5)^2*pi^2(0.88)=1.409684e+00
    "000000001011010101",  -- (p-0.5)^2*pi^2(0.88)=1.416979e+00
    "000000001011011001",  -- (p-0.5)^2*pi^2(0.88)=1.424292e+00
    "000000001011011101",  -- (p-0.5)^2*pi^2(0.88)=1.431624e+00
    "000000001011100001",  -- (p-0.5)^2*pi^2(0.88)=1.438975e+00
    "000000001011100101",  -- (p-0.5)^2*pi^2(0.88)=1.446345e+00
    "000000001011101000",  -- (p-0.5)^2*pi^2(0.88)=1.453734e+00
    "000000001011101100",  -- (p-0.5)^2*pi^2(0.88)=1.461141e+00
    "000000001011110000",  -- (p-0.5)^2*pi^2(0.89)=1.468568e+00
    "000000001011110100",  -- (p-0.5)^2*pi^2(0.89)=1.476013e+00
    "000000001011111000",  -- (p-0.5)^2*pi^2(0.89)=1.483477e+00
    "000000001011111011",  -- (p-0.5)^2*pi^2(0.89)=1.490960e+00
    "000000001011111111",  -- (p-0.5)^2*pi^2(0.89)=1.498462e+00
    "000000001100000011",  -- (p-0.5)^2*pi^2(0.89)=1.505982e+00
    "000000001100000111",  -- (p-0.5)^2*pi^2(0.89)=1.513521e+00
    "000000001100001011",  -- (p-0.5)^2*pi^2(0.89)=1.521080e+00
    "000000001100001111",  -- (p-0.5)^2*pi^2(0.89)=1.528657e+00
    "000000001100010011",  -- (p-0.5)^2*pi^2(0.89)=1.536252e+00
    "000000001100010110",  -- (p-0.5)^2*pi^2(0.90)=1.543867e+00
    "000000001100011010",  -- (p-0.5)^2*pi^2(0.90)=1.551500e+00
    "000000001100011110",  -- (p-0.5)^2*pi^2(0.90)=1.559153e+00
    "000000001100100010",  -- (p-0.5)^2*pi^2(0.90)=1.566824e+00
    "000000001100100110",  -- (p-0.5)^2*pi^2(0.90)=1.574514e+00
    "000000001100101010",  -- (p-0.5)^2*pi^2(0.90)=1.582222e+00
    "000000001100101110",  -- (p-0.5)^2*pi^2(0.90)=1.589950e+00
    "000000001100110010",  -- (p-0.5)^2*pi^2(0.90)=1.597696e+00
    "000000001100110110",  -- (p-0.5)^2*pi^2(0.90)=1.605462e+00
    "000000001100111010",  -- (p-0.5)^2*pi^2(0.90)=1.613246e+00
    "000000001100111110",  -- (p-0.5)^2*pi^2(0.91)=1.621049e+00
    "000000001101000010",  -- (p-0.5)^2*pi^2(0.91)=1.628870e+00
    "000000001101000110",  -- (p-0.5)^2*pi^2(0.91)=1.636711e+00
    "000000001101001010",  -- (p-0.5)^2*pi^2(0.91)=1.644570e+00
    "000000001101001110",  -- (p-0.5)^2*pi^2(0.91)=1.652448e+00
    "000000001101010010",  -- (p-0.5)^2*pi^2(0.91)=1.660345e+00
    "000000001101010110",  -- (p-0.5)^2*pi^2(0.91)=1.668261e+00
    "000000001101011010",  -- (p-0.5)^2*pi^2(0.91)=1.676196e+00
    "000000001101011110",  -- (p-0.5)^2*pi^2(0.91)=1.684149e+00
    "000000001101100010",  -- (p-0.5)^2*pi^2(0.91)=1.692122e+00
    "000000001101100110",  -- (p-0.5)^2*pi^2(0.92)=1.700113e+00
    "000000001101101011",  -- (p-0.5)^2*pi^2(0.92)=1.708123e+00
    "000000001101101111",  -- (p-0.5)^2*pi^2(0.92)=1.716151e+00
    "000000001101110011",  -- (p-0.5)^2*pi^2(0.92)=1.724199e+00
    "000000001101110111",  -- (p-0.5)^2*pi^2(0.92)=1.732265e+00
    "000000001101111011",  -- (p-0.5)^2*pi^2(0.92)=1.740351e+00
    "000000001101111111",  -- (p-0.5)^2*pi^2(0.92)=1.748455e+00
    "000000001110000011",  -- (p-0.5)^2*pi^2(0.92)=1.756578e+00
    "000000001110001000",  -- (p-0.5)^2*pi^2(0.92)=1.764719e+00
    "000000001110001100",  -- (p-0.5)^2*pi^2(0.92)=1.772880e+00
    "000000001110010000",  -- (p-0.5)^2*pi^2(0.92)=1.781059e+00
    "000000001110010100",  -- (p-0.5)^2*pi^2(0.93)=1.789257e+00
    "000000001110011000",  -- (p-0.5)^2*pi^2(0.93)=1.797474e+00
    "000000001110011101",  -- (p-0.5)^2*pi^2(0.93)=1.805710e+00
    "000000001110100001",  -- (p-0.5)^2*pi^2(0.93)=1.813965e+00
    "000000001110100101",  -- (p-0.5)^2*pi^2(0.93)=1.822238e+00
    "000000001110101001",  -- (p-0.5)^2*pi^2(0.93)=1.830531e+00
    "000000001110101101",  -- (p-0.5)^2*pi^2(0.93)=1.838842e+00
    "000000001110110010",  -- (p-0.5)^2*pi^2(0.93)=1.847172e+00
    "000000001110110110",  -- (p-0.5)^2*pi^2(0.93)=1.855521e+00
    "000000001110111010",  -- (p-0.5)^2*pi^2(0.93)=1.863888e+00
    "000000001110111111",  -- (p-0.5)^2*pi^2(0.94)=1.872275e+00
    "000000001111000011",  -- (p-0.5)^2*pi^2(0.94)=1.880680e+00
    "000000001111000111",  -- (p-0.5)^2*pi^2(0.94)=1.889104e+00
    "000000001111001100",  -- (p-0.5)^2*pi^2(0.94)=1.897547e+00
    "000000001111010000",  -- (p-0.5)^2*pi^2(0.94)=1.906009e+00
    "000000001111010100",  -- (p-0.5)^2*pi^2(0.94)=1.914489e+00
    "000000001111011001",  -- (p-0.5)^2*pi^2(0.94)=1.922989e+00
    "000000001111011101",  -- (p-0.5)^2*pi^2(0.94)=1.931507e+00
    "000000001111100001",  -- (p-0.5)^2*pi^2(0.94)=1.940044e+00
    "000000001111100110",  -- (p-0.5)^2*pi^2(0.94)=1.948600e+00
    "000000001111101010",  -- (p-0.5)^2*pi^2(0.95)=1.957174e+00
    "000000001111101110",  -- (p-0.5)^2*pi^2(0.95)=1.965768e+00
    "000000001111110011",  -- (p-0.5)^2*pi^2(0.95)=1.974380e+00
    "000000001111110111",  -- (p-0.5)^2*pi^2(0.95)=1.983011e+00
    "000000001111111100",  -- (p-0.5)^2*pi^2(0.95)=1.991661e+00
    "000000010000000000",  -- (p-0.5)^2*pi^2(0.95)=2.000330e+00
    "000000010000000101",  -- (p-0.5)^2*pi^2(0.95)=2.009018e+00
    "000000010000001001",  -- (p-0.5)^2*pi^2(0.95)=2.017724e+00
    "000000010000001110",  -- (p-0.5)^2*pi^2(0.95)=2.026450e+00
    "000000010000010010",  -- (p-0.5)^2*pi^2(0.95)=2.035194e+00
    "000000010000010111",  -- (p-0.5)^2*pi^2(0.96)=2.043957e+00
    "000000010000011011",  -- (p-0.5)^2*pi^2(0.96)=2.052738e+00
    "000000010000100000",  -- (p-0.5)^2*pi^2(0.96)=2.061539e+00
    "000000010000100100",  -- (p-0.5)^2*pi^2(0.96)=2.070358e+00
    "000000010000101001",  -- (p-0.5)^2*pi^2(0.96)=2.079197e+00
    "000000010000101101",  -- (p-0.5)^2*pi^2(0.96)=2.088054e+00
    "000000010000110010",  -- (p-0.5)^2*pi^2(0.96)=2.096929e+00
    "000000010000110110",  -- (p-0.5)^2*pi^2(0.96)=2.105824e+00
    "000000010000111011",  -- (p-0.5)^2*pi^2(0.96)=2.114738e+00
    "000000010000111111",  -- (p-0.5)^2*pi^2(0.96)=2.123670e+00
    "000000010001000100",  -- (p-0.5)^2*pi^2(0.96)=2.132621e+00
    "000000010001001000",  -- (p-0.5)^2*pi^2(0.97)=2.141591e+00
    "000000010001001101",  -- (p-0.5)^2*pi^2(0.97)=2.150580e+00
    "000000010001010010",  -- (p-0.5)^2*pi^2(0.97)=2.159588e+00
    "000000010001010110",  -- (p-0.5)^2*pi^2(0.97)=2.168614e+00
    "000000010001011011",  -- (p-0.5)^2*pi^2(0.97)=2.177660e+00
    "000000010001100000",  -- (p-0.5)^2*pi^2(0.97)=2.186724e+00
    "000000010001100100",  -- (p-0.5)^2*pi^2(0.97)=2.195807e+00
    "000000010001101001",  -- (p-0.5)^2*pi^2(0.97)=2.204908e+00
    "000000010001101110",  -- (p-0.5)^2*pi^2(0.97)=2.214029e+00
    "000000010001110010",  -- (p-0.5)^2*pi^2(0.97)=2.223168e+00
    "000000010001110111",  -- (p-0.5)^2*pi^2(0.98)=2.232327e+00
    "000000010001111100",  -- (p-0.5)^2*pi^2(0.98)=2.241504e+00
    "000000010010000000",  -- (p-0.5)^2*pi^2(0.98)=2.250700e+00
    "000000010010000101",  -- (p-0.5)^2*pi^2(0.98)=2.259914e+00
    "000000010010001010",  -- (p-0.5)^2*pi^2(0.98)=2.269148e+00
    "000000010010001111",  -- (p-0.5)^2*pi^2(0.98)=2.278400e+00
    "000000010010010011",  -- (p-0.5)^2*pi^2(0.98)=2.287672e+00
    "000000010010011000",  -- (p-0.5)^2*pi^2(0.98)=2.296962e+00
    "000000010010011101",  -- (p-0.5)^2*pi^2(0.98)=2.306270e+00
    "000000010010100010",  -- (p-0.5)^2*pi^2(0.98)=2.315598e+00
    "000000010010100110",  -- (p-0.5)^2*pi^2(0.99)=2.324945e+00
    "000000010010101011",  -- (p-0.5)^2*pi^2(0.99)=2.334310e+00
    "000000010010110000",  -- (p-0.5)^2*pi^2(0.99)=2.343694e+00
    "000000010010110101",  -- (p-0.5)^2*pi^2(0.99)=2.353097e+00
    "000000010010111010",  -- (p-0.5)^2*pi^2(0.99)=2.362519e+00
    "000000010010111110",  -- (p-0.5)^2*pi^2(0.99)=2.371959e+00
    "000000010011000011",  -- (p-0.5)^2*pi^2(0.99)=2.381419e+00
    "000000010011001000",  -- (p-0.5)^2*pi^2(0.99)=2.390897e+00
    "000000010011001101",  -- (p-0.5)^2*pi^2(0.99)=2.400394e+00
    "000000010011010010",  -- (p-0.5)^2*pi^2(0.99)=2.409910e+00
    "000000010011010111",  -- (p-0.5)^2*pi^2(1.00)=2.419445e+00
    "000000010011011100",  -- (p-0.5)^2*pi^2(1.00)=2.428999e+00
    "000000010011100001",  -- (p-0.5)^2*pi^2(1.00)=2.438571e+00
    "000000010011100101",  -- (p-0.5)^2*pi^2(1.00)=2.448162e+00
    "000000010011101010"   -- (p-0.5)^2*pi^2(1.00)=2.457772e+00
    );

  constant CI_ROM_INIT : t_BRAM18k_init_val := fn_BRAM18k_conv_10_18_to_init(
    p_10_18_init_val => ci_data_table
    );
begin

  NON_ZERO_LAT : if (C_LATENCY /= 0) generate
    -- purpose : force model to be RTL on spartan3, as problems wit xbip_bram18k
    function fn_get_model_type(p_model_type : integer; p_xdf : string) return integer is
      variable model_type : integer;
    begin
      if derived(p_xdf, "spartan3") then
        model_type := 1;  -- RTL
      else
        model_type := p_model_type;
      end if;
      return model_type;
    end function fn_get_model_type;

    constant CI_LOC_MODEL_TYPE  : integer := fn_get_model_type(C_MODEL_TYPE, C_XDEVICEFAMILY);
    constant CI_SUPPORTS_DSP48A : boolean := supports_dsp48a(C_XDEVICEFAMILY)>1; 
    constant CI_RTL             : boolean := derived(C_XDEVICEFAMILY, "spartan3") or CI_SUPPORTS_DSP48A;
  begin
    RTL_ROM : if CI_RTL generate
      L1 : if C_LATENCY = 1 generate
        OP_REG : process (CLK)
       begin
         if rising_edge(CLK) then
          if CE='1' then
              D  <= ci_data_table(to_integer(unsigned(A)));
          end if;
        end if;
       end process OP_REG;
     end generate L1;

     L2 : if C_LATENCY >= 2 generate
       signal data1  : std_logic_vector(17 downto 0);  
        signal data2  : std_logic_vector(17 downto 0);  
     begin
   
       OP1_REG : process (CLK)
       begin
         if rising_edge(CLK) then
           if CE='1' then
             data1  <= ci_data_table(to_integer(unsigned(A)));
           end if;
         end if;
       end process OP1_REG;

       OP2_REG : process (CLK)
       begin
         if rising_edge(CLK) then
          if CE='1' then
            data2 <= data1;
          end if;
        end if;
       end process OP2_REG;

       EXTRA_REG : xbip_pipe_v2_0_xst
         generic map(
           C_LATENCY  => C_LATENCY-2,
           C_HAS_CE   => 1,
           C_WIDTH    => 18
         )
         port map(
           CLK  => CLK,
           CE   => CE,
           D    => data2,
           Q    => D
         );
     end generate L2;
   end generate RTL_ROM;
   
   STRUCT_ROM : if not(CI_RTL) generate
     I_BROM : xbip_bram18k_v2_1_xst
       generic map(
         C_XDEVICEFAMILY => C_XDEVICEFAMILY,
         C_VERBOSITY     => 0,
         C_OPTIMIZE_GOAL => 0,
         C_MODEL_TYPE    => CI_LOC_MODEL_TYPE,
         C_LATENCY       => C_LATENCY,
         C_ADDR_WIDTH    => 10,
         C_DATA_WIDTH    => 18,
         C_INIT_VAL      => CI_ROM_INIT
         )
       port map(
         CLK      => CLK,
         CE       => CE,
         SCLR     => SCLR,
         ADDR1    => A,
         DATAOUT1 => D
         );
    end generate STRUCT_ROM;
  end generate NON_ZERO_LAT;

  ZERO_LAT: if C_LATENCY = 0 generate
    signal AI : integer range 0 to 1023 := 0;
  begin

    AI <= to_integer(unsigned(A));
    D  <= ci_data_table(AI);

  end generate ZERO_LAT;
end rtl;
