// --------------------------------------------------------------------
// >>>>>>>>>>>>>>>>>>>>>>>>> COPYRIGHT NOTICE <<<<<<<<<<<<<<<<<<<<<<<<<
// --------------------------------------------------------------------
// Copyright (c) 2005 by Lattice Semiconductor Corporation
// --------------------------------------------------------------------
//
//
//                     Lattice Semiconductor Corporation
//                     5555 NE Moore Court
//                     Hillsboro, OR 97214
//                     U.S.A.
//
//                     TEL: 1-800-Lattice  (USA and Canada)
//                          1-408-826-6000 (other locations)
//
//                     web: http://www.latticesemi.com/
//                     email: techsupport@latticesemi.com
//
// --------------------------------------------------------------------
//
// Simulation Library File for ORCA4
//
// $Header: /home/dmsys/pvcs/RCSMigTest/rcs/verilog/pkg/versclibs/data/orca4/RCS/ULIS.v,v 1.2 2005/05/19 19:02:19 pradeep Exp $ 
//
`timescale 1 ns / 1 ps

`celldefine

module ULIS (RDATA0, RDATA1, RDATA2, RDATA3, RDATA4, RDATA5, RDATA6, RDATA7, RDATA8,
             RDATA9, RDATA10, RDATA11, RDATA12, RDATA13, RDATA14, RDATA15, RDATA16, RDATA17,
             RDATA18, RDATA19, RDATA20, RDATA21, RDATA22, RDATA23, RDATA24, RDATA25,
             RDATA26, RDATA27, RDATA28, RDATA29, RDATA30, RDATA31, RDATA32, RDATA33,
             RDATA34, RDATA35, CLK, RESET, ACK, RETRY, ERR, IRQ, SWDATA0, SWDATA1, SWDATA2,
             SWDATA3, SWDATA4, SWDATA5, SWDATA6, SWDATA7, SWDATA8, SWDATA9, SWDATA10, 
             SWDATA11, SWDATA12, SWDATA13, SWDATA14, SWDATA15, SWDATA16, SWDATA17, SWDATA18,
             SWDATA19, SWDATA20, SWDATA21, SWDATA22, SWDATA23, SWDATA24, SWDATA25,
             SWDATA26, SWDATA27, SWDATA28, SWDATA29, SWDATA30, SWDATA31, SWDATA32, SWDATA33,
             SWDATA34, SWDATA35, SADDR0, SADDR1, SADDR2, SADDR3, SADDR4, SADDR5, SADDR6,
             SADDR7, SADDR8, SADDR9, SADDR10, SADDR11, SADDR12, SADDR13, SADDR14, SADDR15,
             SADDR16, SADDR17, SBURST, SRDY, SWR, SSIZE0, SSIZE1,
             WDATA0, WDATA1, WDATA2, WDATA3, WDATA4, WDATA5, WDATA6, WDATA7, WDATA8,
             WDATA9, WDATA10, WDATA11, WDATA12, WDATA13, WDATA14, WDATA15, WDATA16, WDATA17,
             WDATA18, WDATA19, WDATA20, WDATA21, WDATA22, WDATA23, WDATA24, WDATA25,
             WDATA26, WDATA27, WDATA28, WDATA29, WDATA30, WDATA31, WDATA32, WDATA33,
             WDATA34, WDATA35, ADDR0, ADDR1, ADDR2, ADDR3, ADDR4, ADDR5, ADDR6, ADDR7,
             ADDR8, ADDR9, ADDR10, ADDR11, ADDR12, ADDR13, ADDR14, ADDR15, ADDR16,
             ADDR17, BURST, RDY, WR, SIZE0, SIZE1, SRDATA0, SRDATA1, SRDATA2, SRDATA3,
             SRDATA4, SRDATA5, SRDATA6, SRDATA7, SRDATA8, SRDATA9, SRDATA10, SRDATA11,
             SRDATA12, SRDATA13, SRDATA14, SRDATA15, SRDATA16, SRDATA17, SRDATA18, SRDATA19,
             SRDATA20, SRDATA21, SRDATA22, SRDATA23, SRDATA24, SRDATA25, SRDATA26, SRDATA27,
             SRDATA28, SRDATA29, SRDATA30, SRDATA31, SRDATA32, SRDATA33, SRDATA34, SRDATA35,
             SCLK, SRESET, SACK, SRETRY, SERR, SIRQ);

input RDATA0, RDATA1, RDATA2, RDATA3, RDATA4, RDATA5, RDATA6, RDATA7, RDATA8;
input RDATA9, RDATA10, RDATA11, RDATA12, RDATA13, RDATA14, RDATA15, RDATA16, RDATA17;
input RDATA18, RDATA19, RDATA20, RDATA21, RDATA22, RDATA23, RDATA24, RDATA25, RDATA26;
input RDATA27, RDATA28, RDATA29, RDATA30, RDATA31, RDATA32, RDATA33, RDATA34, RDATA35;
input CLK, RESET, ACK, RETRY, ERR, IRQ, SWDATA0, SWDATA1, SWDATA2, SWDATA3, SWDATA4;
input SWDATA5, SWDATA6, SWDATA7, SWDATA8, SWDATA9, SWDATA10, SWDATA11, SWDATA12;
input SWDATA13, SWDATA14, SWDATA15, SWDATA16, SWDATA17, SWDATA18, SWDATA19, SWDATA20;
input SWDATA21, SWDATA22, SWDATA23, SWDATA24, SWDATA25, SWDATA26, SWDATA27, SWDATA28;
input SWDATA29, SWDATA30, SWDATA31, SWDATA32, SWDATA33, SWDATA34, SWDATA35, SADDR0;
input SADDR1, SADDR2, SADDR3, SADDR4, SADDR5, SADDR6, SADDR7, SADDR8, SADDR9, SADDR10;
input SADDR11, SADDR12, SADDR13, SADDR14, SADDR15, SADDR16, SADDR17, SBURST;
input SRDY, SWR, SSIZE0, SSIZE1;

output WDATA0, WDATA1, WDATA2, WDATA3, WDATA4, WDATA5, WDATA6, WDATA7, WDATA8, WDATA9;
output WDATA10, WDATA11, WDATA12, WDATA13, WDATA14, WDATA15, WDATA16, WDATA17, WDATA18;
output WDATA19, WDATA20, WDATA21, WDATA22, WDATA23, WDATA24, WDATA25, WDATA26, WDATA27;
output WDATA28, WDATA29, WDATA30, WDATA31, WDATA32, WDATA33, WDATA34, WDATA35;
output ADDR0, ADDR1, ADDR2, ADDR3, ADDR4, ADDR5, ADDR6, ADDR7, ADDR8, ADDR9;
output ADDR10, ADDR11, ADDR12, ADDR13, ADDR14, ADDR15, ADDR16, ADDR17, BURST, RDY;
output WR, SIZE0, SIZE1, SRDATA0, SRDATA1, SRDATA2, SRDATA3, SRDATA4, SRDATA5;
output SRDATA6, SRDATA7, SRDATA8, SRDATA9, SRDATA10, SRDATA11, SRDATA12, SRDATA13, SRDATA14;
output SRDATA15, SRDATA16, SRDATA17, SRDATA18, SRDATA19, SRDATA20, SRDATA21, SRDATA22;
output SRDATA23, SRDATA24, SRDATA25, SRDATA26, SRDATA27, SRDATA28, SRDATA29, SRDATA30;
output SRDATA31, SRDATA32, SRDATA33, SRDATA34, SRDATA35, SCLK, SRESET;
output SACK, SRETRY, SERR, SIRQ;

  buf  (WDATA0, SWDATA0);
  buf  (WDATA1, SWDATA1);
  buf  (WDATA2, SWDATA2);
  buf  (WDATA3, SWDATA3);
  buf  (WDATA4, SWDATA4);
  buf  (WDATA5, SWDATA5);
  buf  (WDATA6, SWDATA6);
  buf  (WDATA7, SWDATA7);
  buf  (WDATA8, SWDATA8);
  buf  (WDATA9, SWDATA9);
  buf  (WDATA10, SWDATA10);
  buf  (WDATA11, SWDATA11);
  buf  (WDATA12, SWDATA12);
  buf  (WDATA13, SWDATA13);
  buf  (WDATA14, SWDATA14);
  buf  (WDATA15, SWDATA15);
  buf  (WDATA16, SWDATA16);
  buf  (WDATA17, SWDATA17);
  buf  (WDATA18, SWDATA18);
  buf  (WDATA19, SWDATA19);
  buf  (WDATA20, SWDATA20);
  buf  (WDATA21, SWDATA21);
  buf  (WDATA22, SWDATA22);
  buf  (WDATA23, SWDATA23);
  buf  (WDATA24, SWDATA24);
  buf  (WDATA25, SWDATA25);
  buf  (WDATA26, SWDATA26);
  buf  (WDATA27, SWDATA27);
  buf  (WDATA28, SWDATA28);
  buf  (WDATA29, SWDATA29);
  buf  (WDATA30, SWDATA30);
  buf  (WDATA31, SWDATA31);
  buf  (WDATA32, SWDATA32);
  buf  (WDATA33, SWDATA33);
  buf  (WDATA34, SWDATA34);
  buf  (WDATA35, SWDATA35);
  buf  (BURST, SBURST);
  buf  (RDY, SRDY);
  buf  (WR, SWR);
  buf  (SIZE0, SSIZE0);
  buf  (SIZE1, SSIZE1);
  buf  (ADDR0, SADDR0);
  buf  (ADDR1, SADDR1);
  buf  (ADDR2, SADDR2);
  buf  (ADDR3, SADDR3);
  buf  (ADDR4, SADDR4);
  buf  (ADDR5, SADDR5);
  buf  (ADDR6, SADDR6);
  buf  (ADDR7, SADDR7);
  buf  (ADDR8, SADDR8);
  buf  (ADDR9, SADDR9);
  buf  (ADDR10, SADDR10);
  buf  (ADDR11, SADDR11);
  buf  (ADDR12, SADDR12);
  buf  (ADDR13, SADDR13);
  buf  (ADDR14, SADDR14);
  buf  (ADDR15, SADDR15);
  buf  (ADDR16, SADDR16);
  buf  (ADDR17, SADDR17);
  buf  (SRDATA0, RDATA0);
  buf  (SRDATA1, RDATA1);
  buf  (SRDATA2, RDATA2);
  buf  (SRDATA3, RDATA3);
  buf  (SRDATA4, RDATA4);
  buf  (SRDATA5, RDATA5);
  buf  (SRDATA6, RDATA6);
  buf  (SRDATA7, RDATA7);
  buf  (SRDATA8, RDATA8);
  buf  (SRDATA9, RDATA9);
  buf  (SRDATA10, RDATA10);
  buf  (SRDATA11, RDATA11);
  buf  (SRDATA12, RDATA12);
  buf  (SRDATA13, RDATA13);
  buf  (SRDATA14, RDATA14);
  buf  (SRDATA15, RDATA15);
  buf  (SRDATA16, RDATA16);
  buf  (SRDATA17, RDATA17);
  buf  (SRDATA18, RDATA18);
  buf  (SRDATA19, RDATA19);
  buf  (SRDATA20, RDATA20);
  buf  (SRDATA21, RDATA21);
  buf  (SRDATA22, RDATA22);
  buf  (SRDATA23, RDATA23);
  buf  (SRDATA24, RDATA24);
  buf  (SRDATA25, RDATA25);
  buf  (SRDATA26, RDATA26);
  buf  (SRDATA27, RDATA27);
  buf  (SRDATA28, RDATA28);
  buf  (SRDATA29, RDATA29);
  buf  (SRDATA30, RDATA30);
  buf  (SRDATA31, RDATA31);
  buf  (SRDATA32, RDATA32);
  buf  (SRDATA33, RDATA33);
  buf  (SRDATA34, RDATA34);
  buf  (SRDATA35, RDATA35);
  buf  (SCLK, CLK);
  buf  (SRESET, RESET);
  buf  (SACK, ACK);
  buf  (SRETRY, RETRY);
  buf  (SERR, ERR);
  buf  (SIRQ, IRQ);

endmodule

`endcelldefine

