*  
* Diode Model Produced by Altium Ltd  
* Date:  3-May-2004 
*  
* Manufacturer: Renesas  
* Component Name: HDSP-7401  
*  
* Parameters derived from information available in data sheet.  
* 
*                 common-anode
*                 |  cathode-f
*                 |  |  cathode-g
*                 |  |  |  cathode-e
*                 |  |  |  |  cathode-d
*                 |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  |  cathode-c
*                 |  |  |  |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_7401 1  2  3  4  5  6  7  8  9  10

DA1  1  10  dHDSP_7401
DB1  1   9  dHDSP_7401
DC1  1   8  dHDSP_7401
DD1  1   5  dHDSP_7401
DE1  1   4  dHDSP_7401
DF1  1   2  dHDSP_7401
DG1  1   3  dHDSP_7401
DDP1 1   7  dHDSP_7401

DA2  6  10  dHDSP_7401
DB2  6   9  dHDSP_7401
DC2  6   8  dHDSP_7401
DD2  6   5  dHDSP_7401
DE2  6   4  dHDSP_7401
DF2  6   2  dHDSP_7401
DG2  6   3  dHDSP_7401
DDP2 6   7  dHDSP_7401

.MODEL dHDSP_7401 D
+ (  
+    IS = 2.77296438E-23 
+    N  = 1.39205436 
+    RS = 25.13253104 
+    BV = 45.00000000 
+    IBV = 100u 
+ )  

.ENDS HDSP_7401