*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-A513  
*  
* Parameters derived from information available in data sheet.  
*
*                 common-cathode
*                 |  anode-f
*                 |  |  anode-g
*                 |  |  |  anode-e
*                 |  |  |  |  anode-d
*                 |  |  |  |  |  common-cathode
*                 |  |  |  |  |  |  anode-DP
*                 |  |  |  |  |  |  |  anode-c
*                 |  |  |  |  |  |  |  |  anode-b
*                 |  |  |  |  |  |  |  |  |  anode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_A513 1  2  3  4  5  6  7  8  9  10

DA1  10  1 dHDSP_A513
DB1   9  1 dHDSP_A513
DC1   8  1 dHDSP_A513
DD1   5  1 dHDSP_A513
DE1   4  1 dHDSP_A513
DF1   2  1 dHDSP_A513
DG1   3  1 dHDSP_A513
DDP1  7  1 dHDSP_A513

DA2  10  6 dHDSP_A513
DB2   9  6 dHDSP_A513
DC2   8  6 dHDSP_A513
DD2   5  6 dHDSP_A513
DE2   4  6 dHDSP_A513
DF2   2  6 dHDSP_A513
DG2   3  6 dHDSP_A513
DDP2  7  6 dHDSP_A513

.MODEL dHDSP_A513 D
+ (  
+     IS = 1.61114016E-27 
+      N = 1.30291189 
+     RS = 12.83456794 
+     BV = 50 
+    IBV = 100u 
+ )   

.ENDS HDSP_A513