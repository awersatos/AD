*Vacuum Tube Dual Triode (Audio freq.)
*Connections:
*              Plate 1
*              | Grid 1
*              | | Cathode 1
*              | | | Plate 2
*              | | | | Grid 2
*              | | | | | Cathode 2
*              | | | | | | H H HM
*              | | | | | | | | |
.SUBCKT 12AU7  1 2 3 6 7 8 4 5 9
X1 1 2 3 12AU7s
X2 6 7 8 12AU7s
RH1 4 9 100
RH2 5 9 100
.ENDS 12AU7

*Vacuum Tube Triode (Audio freq.)
*Connections:
*              Plate
*              | Grid
*              | | Cathode
*              | | |
.SUBCKT 12AU7s 1 3 4
B1 2 4 I=((URAMP((V(2,4)/18)+V(3,4)))^1.5)/1151
C1 3 4 1.6E-12
C2 3 1 1.5E-12
C3 1 4 0.5E-12
R1 3 5 10E+3
D1 1 2 DX
D2 4 2 DX2
D3 5 4 DX
.MODEL DX D(IS=1.0E-12 RS=1.0)
.MODEL DX2 D(IS=1.0E-9 RS=1.0)
.ENDS 12AU7s
