*  
* Diode Model Produced by Altium Ltd  
* Date:  10-Mar-2004 
*  
* Manufacturer: Agilent  
* Component Name: HDSP-A211  
*  
* Parameters derived from information available in data sheet.  
*
*                 common-anode
*                 |  cathode-f
*                 |  |  cathode-g
*                 |  |  |  cathode-e
*                 |  |  |  |  cathode-d
*                 |  |  |  |  |  common-anode
*                 |  |  |  |  |  |  cathode-DP
*                 |  |  |  |  |  |  |  cathode-c
*                 |  |  |  |  |  |  |  |  cathode-b
*                 |  |  |  |  |  |  |  |  |  cathode-a
*                 |  |  |  |  |  |  |  |  |  |
.SUBCKT HDSP_A211 1  2  3  4  5  6  7  8  9  10

DA1  1  10 dHDSP_A211
DB1  1   9 dHDSP_A211
DC1  1   8 dHDSP_A211
DD1  1   5 dHDSP_A211
DE1  1   4 dHDSP_A211
DF1  1   2 dHDSP_A211
DG1  1   3 dHDSP_A211
DDP1 1   7 dHDSP_A211

DA2  6  10 dHDSP_A211
DB2  6   9 dHDSP_A211
DC2  6   8 dHDSP_A211
DD2  6   5 dHDSP_A211
DE2  6   4 dHDSP_A211
DF2  6   2 dHDSP_A211
DG2  6   3 dHDSP_A211
DDP2 6   7 dHDSP_A211

.MODEL dHDSP_A211 D
+ (  
+     IS = 2.92097419E-52 
+      N = 0.52799867 
+     RS = 25.27044243 
+     BV = 30
+    IBV = 100u 
+ )  

.ENDS HDSP_A211