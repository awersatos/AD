-------------------------------------------------------
--  Copyright (c) 1995/2006 Xilinx Inc.
--  All Right Reserved.
-------------------------------------------------------
--
--   ____  ____
--  /   /\/   / 
-- /___/  \  /     Vendor      : Xilinx 
-- \   \   \/      Version : 11.1
--  \   \          Description : 
--  /   /                      
-- /___/   /\      Filename    : X_PPC440.vhd
-- \   \  /  \     Timestamp   : Fri Apr 20 15:15:22 2007

--  \__ \/\__ \                   
--                                 
--  Generated by    : write_vhdl
--  Revision: 
-------------------------------------------------------

----- CELL X_PPC440 -----

library IEEE;
use IEEE.STD_LOGIC_1164.all;

library IEEE;
use IEEE.VITAL_Timing.all;

library simprim;
use simprim.VCOMPONENTS.all; 

library secureip; 
use secureip.all; 

entity X_PPC440 is
generic (
	TimingChecksOn : boolean := TRUE;
	InstancePath   : string  := "*";
	Xon            : boolean := TRUE;
	MsgOn          : boolean := FALSE;

	LOC             : string  := "UNPLACED";

	APU_CONTROL : bit_vector := X"02000";
	APU_UDI0 : bit_vector := X"000000";
	APU_UDI1 : bit_vector := X"000000";
	APU_UDI10 : bit_vector := X"000000";
	APU_UDI11 : bit_vector := X"000000";
	APU_UDI12 : bit_vector := X"000000";
	APU_UDI13 : bit_vector := X"000000";
	APU_UDI14 : bit_vector := X"000000";
	APU_UDI15 : bit_vector := X"000000";
	APU_UDI2 : bit_vector := X"000000";
	APU_UDI3 : bit_vector := X"000000";
	APU_UDI4 : bit_vector := X"000000";
	APU_UDI5 : bit_vector := X"000000";
	APU_UDI6 : bit_vector := X"000000";
	APU_UDI7 : bit_vector := X"000000";
	APU_UDI8 : bit_vector := X"000000";
	APU_UDI9 : bit_vector := X"000000";
	CLOCK_DELAY : boolean := FALSE;
	DCR_AUTOLOCK_ENABLE : boolean := TRUE;
	DMA0_CONTROL : bit_vector := X"00";
	DMA0_RXCHANNELCTRL : bit_vector := X"01010000";
	DMA0_RXIRQTIMER : bit_vector := X"3FF";
	DMA0_TXCHANNELCTRL : bit_vector := X"01010000";
	DMA0_TXIRQTIMER : bit_vector := X"3FF";
	DMA1_CONTROL : bit_vector := X"00";
	DMA1_RXCHANNELCTRL : bit_vector := X"01010000";
	DMA1_RXIRQTIMER : bit_vector := X"3FF";
	DMA1_TXCHANNELCTRL : bit_vector := X"01010000";
	DMA1_TXIRQTIMER : bit_vector := X"3FF";
	DMA2_CONTROL : bit_vector := X"00";
	DMA2_RXCHANNELCTRL : bit_vector := X"01010000";
	DMA2_RXIRQTIMER : bit_vector := X"3FF";
	DMA2_TXCHANNELCTRL : bit_vector := X"01010000";
	DMA2_TXIRQTIMER : bit_vector := X"3FF";
	DMA3_CONTROL : bit_vector := X"00";
	DMA3_RXCHANNELCTRL : bit_vector := X"01010000";
	DMA3_RXIRQTIMER : bit_vector := X"3FF";
	DMA3_TXCHANNELCTRL : bit_vector := X"01010000";
	DMA3_TXIRQTIMER : bit_vector := X"3FF";
	INTERCONNECT_IMASK : bit_vector := X"FFFFFFFF";
	INTERCONNECT_TMPL_SEL : bit_vector := X"3FFFFFFF";
	MI_ARBCONFIG : bit_vector := X"00432010";
	MI_BANKCONFLICT_MASK : bit_vector := X"00000000";
	MI_CONTROL : bit_vector := X"0000008F";
	MI_ROWCONFLICT_MASK : bit_vector := X"00000000";
	PPCDM_ASYNCMODE : boolean := FALSE;
	PPCDS_ASYNCMODE : boolean := FALSE;
	PPCM_ARBCONFIG : bit_vector := X"00432010";
	PPCM_CONTROL : bit_vector := X"8000009F";
	PPCM_COUNTER : bit_vector := X"00000500";
	PPCS0_ADDRMAP_TMPL0 : bit_vector := X"FFFFFFFF";
	PPCS0_ADDRMAP_TMPL1 : bit_vector := X"FFFFFFFF";
	PPCS0_ADDRMAP_TMPL2 : bit_vector := X"FFFFFFFF";
	PPCS0_ADDRMAP_TMPL3 : bit_vector := X"FFFFFFFF";
	PPCS0_CONTROL : bit_vector := X"8033336C";
	PPCS0_WIDTH_128N64 : boolean := TRUE;
	PPCS1_ADDRMAP_TMPL0 : bit_vector := X"FFFFFFFF";
	PPCS1_ADDRMAP_TMPL1 : bit_vector := X"FFFFFFFF";
	PPCS1_ADDRMAP_TMPL2 : bit_vector := X"FFFFFFFF";
	PPCS1_ADDRMAP_TMPL3 : bit_vector := X"FFFFFFFF";
	PPCS1_CONTROL : bit_vector := X"8033336C";
	PPCS1_WIDTH_128N64 : boolean := TRUE;
	XBAR_ADDRMAP_TMPL0 : bit_vector := X"FFFF0000";
	XBAR_ADDRMAP_TMPL1 : bit_vector := X"00000000";
	XBAR_ADDRMAP_TMPL2 : bit_vector := X"00000000";
	XBAR_ADDRMAP_TMPL3 : bit_vector := X"00000000";

	tperiod_CPMC440TIMERCLOCK_posedge : VitalDelayType := 0 ps;
	tperiod_CPMDCRCLK_posedge : VitalDelayType := 0 ps;
	tperiod_CPMFCMCLK_posedge : VitalDelayType := 0 ps;
	tperiod_CPMINTERCONNECTCLK_posedge : VitalDelayType := 0 ps;
	tperiod_CPMMCCLK_posedge : VitalDelayType := 0 ps;
	tperiod_CPMPPCMPLBCLK_posedge : VitalDelayType := 0 ps;
	tperiod_CPMPPCS0PLBCLK_posedge : VitalDelayType := 0 ps;
	tperiod_CPMPPCS1PLBCLK_posedge : VitalDelayType := 0 ps;

	tipd_CPMC440CLK : VitalDelayType01 :=  (0 ps, 0 ps);
	tipd_CPMC440CLKEN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_CPMC440CORECLOCKINACTIVE : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_CPMC440TIMERCLOCK : VitalDelayType01 :=  (0 ps, 0 ps);
	tipd_CPMDCRCLK : VitalDelayType01 :=  (0 ps, 0 ps);
	tipd_CPMDMA0LLCLK : VitalDelayType01 :=  (0 ps, 0 ps);
	tipd_CPMDMA1LLCLK : VitalDelayType01 :=  (0 ps, 0 ps);
	tipd_CPMDMA2LLCLK : VitalDelayType01 :=  (0 ps, 0 ps);
	tipd_CPMDMA3LLCLK : VitalDelayType01 :=  (0 ps, 0 ps);
	tipd_CPMFCMCLK : VitalDelayType01 :=  (0 ps, 0 ps);
	tipd_CPMINTERCONNECTCLK : VitalDelayType01 :=  (0 ps, 0 ps);
	tipd_CPMINTERCONNECTCLKEN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_CPMINTERCONNECTCLKNTO1 : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_CPMMCCLK : VitalDelayType01 :=  (0 ps, 0 ps);
	tipd_CPMPPCMPLBCLK : VitalDelayType01 :=  (0 ps, 0 ps);
	tipd_CPMPPCS0PLBCLK : VitalDelayType01 :=  (0 ps, 0 ps);
	tipd_CPMPPCS1PLBCLK : VitalDelayType01 :=  (0 ps, 0 ps);
	tipd_DBGC440DEBUGHALT : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_DBGC440SYSTEMSTATUS : VitalDelayArrayType01 (0 to 4) := (others => (100 ps, 100 ps));
	tipd_DBGC440UNCONDDEBUGEVENT : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_DCRPPCDMACK : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_DCRPPCDMDBUSIN : VitalDelayArrayType01 (0 to 31) := (others => (100 ps, 100 ps));
	tipd_DCRPPCDMTIMEOUTWAIT : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_DCRPPCDSABUS : VitalDelayArrayType01 (0 to 9) := (others => (100 ps, 100 ps));
	tipd_DCRPPCDSDBUSOUT : VitalDelayArrayType01 (0 to 31) := (others => (100 ps, 100 ps));
	tipd_DCRPPCDSREAD : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_DCRPPCDSWRITE : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_EICC440CRITIRQ : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_EICC440EXTIRQ : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_FCMAPUCONFIRMINSTR : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_FCMAPUCR : VitalDelayArrayType01 (0 to 3) := (others => (100 ps, 100 ps));
	tipd_FCMAPUDONE : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_FCMAPUEXCEPTION : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_FCMAPUFPSCRFEX : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_FCMAPURESULT : VitalDelayArrayType01 (0 to 31) := (others => (100 ps, 100 ps));
	tipd_FCMAPURESULTVALID : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_FCMAPUSLEEPNOTREADY : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_FCMAPUSTOREDATA : VitalDelayArrayType01 (0 to 127) := (others => (100 ps, 100 ps));
	tipd_JTGC440TCK : VitalDelayType01 :=  (0 ps, 0 ps);
	tipd_JTGC440TDI : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_JTGC440TMS : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_JTGC440TRSTNEG : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA0RSTENGINEREQ : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA0RXD : VitalDelayArrayType01 (0 to 31) := (others => (100 ps, 100 ps));
	tipd_LLDMA0RXEOFN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA0RXEOPN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA0RXREM : VitalDelayArrayType01 (0 to 3) := (others => (100 ps, 100 ps));
	tipd_LLDMA0RXSOFN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA0RXSOPN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA0RXSRCRDYN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA0TXDSTRDYN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA1RSTENGINEREQ : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA1RXD : VitalDelayArrayType01 (0 to 31) := (others => (100 ps, 100 ps));
	tipd_LLDMA1RXEOFN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA1RXEOPN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA1RXREM : VitalDelayArrayType01 (0 to 3) := (others => (100 ps, 100 ps));
	tipd_LLDMA1RXSOFN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA1RXSOPN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA1RXSRCRDYN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA1TXDSTRDYN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA2RSTENGINEREQ : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA2RXD : VitalDelayArrayType01 (0 to 31) := (others => (100 ps, 100 ps));
	tipd_LLDMA2RXEOFN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA2RXEOPN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA2RXREM : VitalDelayArrayType01 (0 to 3) := (others => (100 ps, 100 ps));
	tipd_LLDMA2RXSOFN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA2RXSOPN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA2RXSRCRDYN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA2TXDSTRDYN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA3RSTENGINEREQ : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA3RXD : VitalDelayArrayType01 (0 to 31) := (others => (100 ps, 100 ps));
	tipd_LLDMA3RXEOFN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA3RXEOPN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA3RXREM : VitalDelayArrayType01 (0 to 3) := (others => (100 ps, 100 ps));
	tipd_LLDMA3RXSOFN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA3RXSOPN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA3RXSRCRDYN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_LLDMA3TXDSTRDYN : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_MCMIADDRREADYTOACCEPT : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_MCMIREADDATA : VitalDelayArrayType01 (0 to 127) := (others => (100 ps, 100 ps));
	tipd_MCMIREADDATAERR : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_MCMIREADDATAVALID : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCMADDRACK : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCMMBUSY : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCMMIRQ : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCMMRDERR : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCMMWRERR : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCMRDBTERM : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCMRDDACK : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCMRDDBUS : VitalDelayArrayType01 (0 to 127) := (others => (100 ps, 100 ps));
	tipd_PLBPPCMRDPENDPRI : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_PLBPPCMRDPENDREQ : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCMRDWDADDR : VitalDelayArrayType01 (0 to 3) := (others => (100 ps, 100 ps));
	tipd_PLBPPCMREARBITRATE : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCMREQPRI : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_PLBPPCMSSIZE : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_PLBPPCMTIMEOUT : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCMWRBTERM : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCMWRDACK : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCMWRPENDPRI : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_PLBPPCMWRPENDREQ : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS0ABORT : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS0ABUS : VitalDelayArrayType01 (0 to 31) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS0BE : VitalDelayArrayType01 (0 to 15) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS0BUSLOCK : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS0LOCKERR : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS0MASTERID : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS0MSIZE : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS0PAVALID : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS0RDBURST : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS0RDPENDPRI : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS0RDPENDREQ : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS0RDPRIM : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS0REQPRI : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS0RNW : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS0SAVALID : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS0SIZE : VitalDelayArrayType01 (0 to 3) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS0TATTRIBUTE : VitalDelayArrayType01 (0 to 15) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS0TYPE : VitalDelayArrayType01 (0 to 2) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS0UABUS : VitalDelayArrayType01 (28 to 31) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS0WRBURST : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS0WRDBUS : VitalDelayArrayType01 (0 to 127) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS0WRPENDPRI : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS0WRPENDREQ : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS0WRPRIM : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS1ABORT : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS1ABUS : VitalDelayArrayType01 (0 to 31) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS1BE : VitalDelayArrayType01 (0 to 15) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS1BUSLOCK : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS1LOCKERR : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS1MASTERID : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS1MSIZE : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS1PAVALID : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS1RDBURST : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS1RDPENDPRI : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS1RDPENDREQ : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS1RDPRIM : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS1REQPRI : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS1RNW : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS1SAVALID : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS1SIZE : VitalDelayArrayType01 (0 to 3) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS1TATTRIBUTE : VitalDelayArrayType01 (0 to 15) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS1TYPE : VitalDelayArrayType01 (0 to 2) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS1UABUS : VitalDelayArrayType01 (28 to 31) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS1WRBURST : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS1WRDBUS : VitalDelayArrayType01 (0 to 127) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS1WRPENDPRI : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_PLBPPCS1WRPENDREQ : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_PLBPPCS1WRPRIM : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_RSTC440RESETCHIP : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_RSTC440RESETCORE : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_RSTC440RESETSYSTEM : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_TIEC440DCURDLDCACHEPLBPRIO : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_TIEC440DCURDNONCACHEPLBPRIO : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_TIEC440DCURDTOUCHPLBPRIO : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_TIEC440DCURDURGENTPLBPRIO : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_TIEC440DCUWRFLUSHPLBPRIO : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_TIEC440DCUWRSTOREPLBPRIO : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_TIEC440DCUWRURGENTPLBPRIO : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_TIEC440ENDIANRESET : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_TIEC440ERPNRESET : VitalDelayArrayType01 (0 to 3) := (others => (100 ps, 100 ps));
	tipd_TIEC440ICURDFETCHPLBPRIO : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_TIEC440ICURDSPECPLBPRIO : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_TIEC440ICURDTOUCHPLBPRIO : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_TIEC440PIR : VitalDelayArrayType01 (28 to 31) := (others => (100 ps, 100 ps));
	tipd_TIEC440PVR : VitalDelayArrayType01 (28 to 31) := (others => (100 ps, 100 ps));
	tipd_TIEC440USERRESET : VitalDelayArrayType01 (0 to 3) := (others => (100 ps, 100 ps));
	tipd_TIEDCRBASEADDR : VitalDelayArrayType01 (0 to 1) := (others => (100 ps, 100 ps));
	tipd_TRCC440TRACEDISABLE : VitalDelayType01 :=  (100 ps, 100 ps);
	tipd_TRCC440TRIGGEREVENTIN : VitalDelayType01 :=  (100 ps, 100 ps);
	tpd_CPMC440CLK_C440CPMCORESLEEPREQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMC440CLK_C440CPMDECIRPTREQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMC440CLK_C440CPMFITIRPTREQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMC440CLK_C440CPMMSRCE : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMC440CLK_C440CPMMSREE : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMC440CLK_C440CPMTIMERRESETREQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMC440CLK_C440CPMWDIRPTREQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMC440CLK_C440DBGSYSTEMCONTROL : VitalDelayArrayType01(0 to 7) := (others => (100 ps, 100 ps));
	tpd_CPMC440CLK_C440MACHINECHECK : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMC440CLK_C440TRCBRANCHSTATUS : VitalDelayArrayType01(0 to 2) := (others => (100 ps, 100 ps));
	tpd_CPMC440CLK_C440TRCCYCLE : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMC440CLK_C440TRCEXECUTIONSTATUS : VitalDelayArrayType01(0 to 4) := (others => (100 ps, 100 ps));
	tpd_CPMC440CLK_C440TRCTRACESTATUS : VitalDelayArrayType01(0 to 6) := (others => (100 ps, 100 ps));
	tpd_CPMC440CLK_C440TRCTRIGGEREVENTOUT : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE : VitalDelayArrayType01(0 to 13) := (others => (100 ps, 100 ps));
	tpd_CPMDCRCLK_PPCDMDCRABUS : VitalDelayArrayType01(0 to 9) := (others => (100 ps, 100 ps));
	tpd_CPMDCRCLK_PPCDMDCRDBUSOUT : VitalDelayArrayType01(0 to 31) := (others => (100 ps, 100 ps));
	tpd_CPMDCRCLK_PPCDMDCRREAD : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDCRCLK_PPCDMDCRUABUS : VitalDelayArrayType01(20 to 21) := (others => (100 ps, 100 ps));
	tpd_CPMDCRCLK_PPCDMDCRWRITE : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDCRCLK_PPCDSDCRACK : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDCRCLK_PPCDSDCRDBUSIN : VitalDelayArrayType01(0 to 31) := (others => (100 ps, 100 ps));
	tpd_CPMDCRCLK_PPCDSDCRTIMEOUTWAIT : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA0LLCLK_DMA0LLRSTENGINEACK : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA0LLCLK_DMA0LLRXDSTRDYN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA0LLCLK_DMA0LLTXD : VitalDelayArrayType01(0 to 31) := (others => (100 ps, 100 ps));
	tpd_CPMDMA0LLCLK_DMA0LLTXEOFN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA0LLCLK_DMA0LLTXEOPN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA0LLCLK_DMA0LLTXREM : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMDMA0LLCLK_DMA0LLTXSOFN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA0LLCLK_DMA0LLTXSOPN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA0LLCLK_DMA0LLTXSRCRDYN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA0LLCLK_DMA0RXIRQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA0LLCLK_DMA0TXIRQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA1LLCLK_DMA1LLRSTENGINEACK : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA1LLCLK_DMA1LLRXDSTRDYN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA1LLCLK_DMA1LLTXD : VitalDelayArrayType01(0 to 31) := (others => (100 ps, 100 ps));
	tpd_CPMDMA1LLCLK_DMA1LLTXEOFN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA1LLCLK_DMA1LLTXEOPN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA1LLCLK_DMA1LLTXREM : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMDMA1LLCLK_DMA1LLTXSOFN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA1LLCLK_DMA1LLTXSOPN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA1LLCLK_DMA1LLTXSRCRDYN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA1LLCLK_DMA1RXIRQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA1LLCLK_DMA1TXIRQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA2LLCLK_DMA2LLRSTENGINEACK : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA2LLCLK_DMA2LLRXDSTRDYN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA2LLCLK_DMA2LLTXD : VitalDelayArrayType01(0 to 31) := (others => (100 ps, 100 ps));
	tpd_CPMDMA2LLCLK_DMA2LLTXEOFN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA2LLCLK_DMA2LLTXEOPN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA2LLCLK_DMA2LLTXREM : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMDMA2LLCLK_DMA2LLTXSOFN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA2LLCLK_DMA2LLTXSOPN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA2LLCLK_DMA2LLTXSRCRDYN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA2LLCLK_DMA2RXIRQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA2LLCLK_DMA2TXIRQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA3LLCLK_DMA3LLRSTENGINEACK : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA3LLCLK_DMA3LLRXDSTRDYN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA3LLCLK_DMA3LLTXD : VitalDelayArrayType01(0 to 31) := (others => (100 ps, 100 ps));
	tpd_CPMDMA3LLCLK_DMA3LLTXEOFN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA3LLCLK_DMA3LLTXEOPN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA3LLCLK_DMA3LLTXREM : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMDMA3LLCLK_DMA3LLTXSOFN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA3LLCLK_DMA3LLTXSOPN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA3LLCLK_DMA3LLTXSRCRDYN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA3LLCLK_DMA3RXIRQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMDMA3LLCLK_DMA3TXIRQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMFCMCLK_APUFCMDECFPUOP : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMFCMCLK_APUFCMDECLDSTXFERSIZE : VitalDelayArrayType01(0 to 2) := (others => (100 ps, 100 ps));
	tpd_CPMFCMCLK_APUFCMDECLOAD : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMFCMCLK_APUFCMDECNONAUTON : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMFCMCLK_APUFCMDECSTORE : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMFCMCLK_APUFCMDECUDI : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMFCMCLK_APUFCMDECUDIVALID : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMFCMCLK_APUFCMENDIAN : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMFCMCLK_APUFCMFLUSH : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMFCMCLK_APUFCMINSTRUCTION : VitalDelayArrayType01(0 to 31) := (others => (100 ps, 100 ps));
	tpd_CPMFCMCLK_APUFCMINSTRVALID : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMFCMCLK_APUFCMLOADBYTEADDR : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMFCMCLK_APUFCMLOADDATA : VitalDelayArrayType01(0 to 127) := (others => (100 ps, 100 ps));
	tpd_CPMFCMCLK_APUFCMLOADDVALID : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMFCMCLK_APUFCMMSRFE0 : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMFCMCLK_APUFCMMSRFE1 : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMFCMCLK_APUFCMNEXTINSTRREADY : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMFCMCLK_APUFCMOPERANDVALID : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMFCMCLK_APUFCMRADATA : VitalDelayArrayType01(0 to 31) := (others => (100 ps, 100 ps));
	tpd_CPMFCMCLK_APUFCMRBDATA : VitalDelayArrayType01(0 to 31) := (others => (100 ps, 100 ps));
	tpd_CPMFCMCLK_APUFCMWRITEBACKOK : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMINTERCONNECTCLK_C440RSTCHIPRESETREQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMINTERCONNECTCLK_C440RSTCORERESETREQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMINTERCONNECTCLK_C440RSTSYSTEMRESETREQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMINTERCONNECTCLK_PPCCPMINTERCONNECTBUSY : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMINTERCONNECTCLK_PPCEICINTERCONNECTIRQ : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMMCCLK_MIMCADDRESS : VitalDelayArrayType01(0 to 35) := (others => (100 ps, 100 ps));
	tpd_CPMMCCLK_MIMCADDRESSVALID : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMMCCLK_MIMCBANKCONFLICT : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMMCCLK_MIMCBYTEENABLE : VitalDelayArrayType01(0 to 15) := (others => (100 ps, 100 ps));
	tpd_CPMMCCLK_MIMCREADNOTWRITE : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMMCCLK_MIMCROWCONFLICT : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMMCCLK_MIMCWRITEDATA : VitalDelayArrayType01(0 to 127) := (others => (100 ps, 100 ps));
	tpd_CPMMCCLK_MIMCWRITEDATAVALID : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCMPLBCLK_PPCMPLBABORT : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCMPLBCLK_PPCMPLBABUS : VitalDelayArrayType01(0 to 31) := (others => (100 ps, 100 ps));
	tpd_CPMPPCMPLBCLK_PPCMPLBBE : VitalDelayArrayType01(0 to 15) := (others => (100 ps, 100 ps));
	tpd_CPMPPCMPLBCLK_PPCMPLBBUSLOCK : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCMPLBCLK_PPCMPLBLOCKERR : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCMPLBCLK_PPCMPLBPRIORITY : VitalDelayArrayType01(0 to 1) := (others => (100 ps, 100 ps));
	tpd_CPMPPCMPLBCLK_PPCMPLBRDBURST : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCMPLBCLK_PPCMPLBREQUEST : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCMPLBCLK_PPCMPLBRNW : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCMPLBCLK_PPCMPLBSIZE : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE : VitalDelayArrayType01(0 to 15) := (others => (100 ps, 100 ps));
	tpd_CPMPPCMPLBCLK_PPCMPLBTYPE : VitalDelayArrayType01(0 to 2) := (others => (100 ps, 100 ps));
	tpd_CPMPPCMPLBCLK_PPCMPLBUABUS : VitalDelayArrayType01(28 to 31) := (others => (100 ps, 100 ps));
	tpd_CPMPPCMPLBCLK_PPCMPLBWRBURST : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS : VitalDelayArrayType01(0 to 127) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS0PLBCLK_PPCS0PLBADDRACK : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS0PLBCLK_PPCS0PLBMBUSY : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS0PLBCLK_PPCS0PLBMIRQ : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS0PLBCLK_PPCS0PLBMRDERR : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS0PLBCLK_PPCS0PLBMWRERR : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS0PLBCLK_PPCS0PLBRDBTERM : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS0PLBCLK_PPCS0PLBRDCOMP : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDACK : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS : VitalDelayArrayType01(0 to 127) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS0PLBCLK_PPCS0PLBRDWDADDR : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS0PLBCLK_PPCS0PLBREARBITRATE : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS0PLBCLK_PPCS0PLBSSIZE : VitalDelayArrayType01(0 to 1) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS0PLBCLK_PPCS0PLBWAIT : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS0PLBCLK_PPCS0PLBWRBTERM : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS0PLBCLK_PPCS0PLBWRCOMP : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS0PLBCLK_PPCS0PLBWRDACK : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS1PLBCLK_PPCS1PLBADDRACK : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS1PLBCLK_PPCS1PLBMBUSY : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS1PLBCLK_PPCS1PLBMIRQ : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS1PLBCLK_PPCS1PLBMRDERR : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS1PLBCLK_PPCS1PLBMWRERR : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS1PLBCLK_PPCS1PLBRDBTERM : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS1PLBCLK_PPCS1PLBRDCOMP : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDACK : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS : VitalDelayArrayType01(0 to 127) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS1PLBCLK_PPCS1PLBRDWDADDR : VitalDelayArrayType01(0 to 3) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS1PLBCLK_PPCS1PLBREARBITRATE : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS1PLBCLK_PPCS1PLBSSIZE : VitalDelayArrayType01(0 to 1) := (others => (100 ps, 100 ps));
	tpd_CPMPPCS1PLBCLK_PPCS1PLBWAIT : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS1PLBCLK_PPCS1PLBWRBTERM : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS1PLBCLK_PPCS1PLBWRCOMP : VitalDelayType01 := (100 ps, 100 ps);
	tpd_CPMPPCS1PLBCLK_PPCS1PLBWRDACK : VitalDelayType01 := (100 ps, 100 ps);
	tpd_JTGC440TCK_C440JTGTDO : VitalDelayType01 := (100 ps, 100 ps);
	tpd_JTGC440TCK_C440JTGTDOEN : VitalDelayType01 := (100 ps, 100 ps);

	thold_CPMC440CORECLOCKINACTIVE_JTGC440TCK_negedge_posedge : VitalDelayType := 0 ps;
	thold_CPMC440CORECLOCKINACTIVE_JTGC440TCK_posedge_posedge : VitalDelayType := 0 ps;
	thold_CPMINTERCONNECTCLKNTO1_CPMINTERCONNECTCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_CPMINTERCONNECTCLKNTO1_CPMINTERCONNECTCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_DBGC440DEBUGHALT_CPMC440CLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_DBGC440DEBUGHALT_CPMC440CLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_DBGC440SYSTEMSTATUS_JTGC440TCK_negedge_posedge : VitalDelayArrayType(0 to 4) := (others => 0 ps);
	thold_DBGC440SYSTEMSTATUS_JTGC440TCK_posedge_posedge : VitalDelayArrayType(0 to 4) := (others => 0 ps);
	thold_DBGC440UNCONDDEBUGEVENT_CPMC440CLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_DBGC440UNCONDDEBUGEVENT_CPMC440CLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_DCRPPCDMACK_CPMDCRCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_DCRPPCDMACK_CPMDCRCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_DCRPPCDMTIMEOUTWAIT_CPMDCRCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_DCRPPCDMTIMEOUTWAIT_CPMDCRCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge : VitalDelayArrayType(0 to 9) := (others => 0 ps);
	thold_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge : VitalDelayArrayType(0 to 9) := (others => 0 ps);
	thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_DCRPPCDSREAD_CPMDCRCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_DCRPPCDSREAD_CPMDCRCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_DCRPPCDSWRITE_CPMDCRCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_DCRPPCDSWRITE_CPMDCRCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_FCMAPUCONFIRMINSTR_CPMFCMCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_FCMAPUCONFIRMINSTR_CPMFCMCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_FCMAPUCR_CPMFCMCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_FCMAPUCR_CPMFCMCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_FCMAPUDONE_CPMFCMCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_FCMAPUDONE_CPMFCMCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_FCMAPUEXCEPTION_CPMFCMCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_FCMAPUEXCEPTION_CPMFCMCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_FCMAPUFPSCRFEX_CPMFCMCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_FCMAPUFPSCRFEX_CPMFCMCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_FCMAPURESULTVALID_CPMFCMCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_FCMAPURESULTVALID_CPMFCMCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_FCMAPUSLEEPNOTREADY_CPMFCMCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_FCMAPUSLEEPNOTREADY_CPMFCMCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	thold_JTGC440TDI_JTGC440TCK_negedge_posedge : VitalDelayType := 0 ps;
	thold_JTGC440TDI_JTGC440TCK_posedge_posedge : VitalDelayType := 0 ps;
	thold_JTGC440TMS_JTGC440TCK_negedge_posedge : VitalDelayType := 0 ps;
	thold_JTGC440TMS_JTGC440TCK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA0RSTENGINEREQ_CPMDMA0LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA0RSTENGINEREQ_CPMDMA0LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_LLDMA0RXEOFN_CPMDMA0LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA0RXEOFN_CPMDMA0LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA0RXEOPN_CPMDMA0LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA0RXEOPN_CPMDMA0LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA0RXREM_CPMDMA0LLCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_LLDMA0RXREM_CPMDMA0LLCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_LLDMA0RXSOFN_CPMDMA0LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA0RXSOFN_CPMDMA0LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA0RXSOPN_CPMDMA0LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA0RXSOPN_CPMDMA0LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA0RXSRCRDYN_CPMDMA0LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA0RXSRCRDYN_CPMDMA0LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA0TXDSTRDYN_CPMDMA0LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA0TXDSTRDYN_CPMDMA0LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA1RSTENGINEREQ_CPMDMA1LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA1RSTENGINEREQ_CPMDMA1LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_LLDMA1RXEOFN_CPMDMA1LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA1RXEOFN_CPMDMA1LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA1RXEOPN_CPMDMA1LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA1RXEOPN_CPMDMA1LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA1RXREM_CPMDMA1LLCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_LLDMA1RXREM_CPMDMA1LLCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_LLDMA1RXSOFN_CPMDMA1LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA1RXSOFN_CPMDMA1LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA1RXSOPN_CPMDMA1LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA1RXSOPN_CPMDMA1LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA1RXSRCRDYN_CPMDMA1LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA1RXSRCRDYN_CPMDMA1LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA1TXDSTRDYN_CPMDMA1LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA1TXDSTRDYN_CPMDMA1LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA2RSTENGINEREQ_CPMDMA2LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA2RSTENGINEREQ_CPMDMA2LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_LLDMA2RXEOFN_CPMDMA2LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA2RXEOFN_CPMDMA2LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA2RXEOPN_CPMDMA2LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA2RXEOPN_CPMDMA2LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA2RXREM_CPMDMA2LLCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_LLDMA2RXREM_CPMDMA2LLCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_LLDMA2RXSOFN_CPMDMA2LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA2RXSOFN_CPMDMA2LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA2RXSOPN_CPMDMA2LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA2RXSOPN_CPMDMA2LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA2RXSRCRDYN_CPMDMA2LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA2RXSRCRDYN_CPMDMA2LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA2TXDSTRDYN_CPMDMA2LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA2TXDSTRDYN_CPMDMA2LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA3RSTENGINEREQ_CPMDMA3LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA3RSTENGINEREQ_CPMDMA3LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_LLDMA3RXEOFN_CPMDMA3LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA3RXEOFN_CPMDMA3LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA3RXEOPN_CPMDMA3LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA3RXEOPN_CPMDMA3LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA3RXREM_CPMDMA3LLCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_LLDMA3RXREM_CPMDMA3LLCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_LLDMA3RXSOFN_CPMDMA3LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA3RXSOFN_CPMDMA3LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA3RXSOPN_CPMDMA3LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA3RXSOPN_CPMDMA3LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA3RXSRCRDYN_CPMDMA3LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA3RXSRCRDYN_CPMDMA3LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA3TXDSTRDYN_CPMDMA3LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_LLDMA3TXDSTRDYN_CPMDMA3LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_MCMIADDRREADYTOACCEPT_CPMMCCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_MCMIADDRREADYTOACCEPT_CPMMCCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_MCMIREADDATAERR_CPMMCCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_MCMIREADDATAERR_CPMMCCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_MCMIREADDATAVALID_CPMMCCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_MCMIREADDATAVALID_CPMMCCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_MCMIREADDATA_CPMMCCLK_negedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	thold_MCMIREADDATA_CPMMCCLK_posedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	thold_PLBPPCMADDRACK_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMADDRACK_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMMBUSY_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMMBUSY_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMMIRQ_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMMIRQ_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMMRDERR_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMMRDERR_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMMWRERR_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMMWRERR_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMRDBTERM_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMRDBTERM_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMRDDACK_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMRDDACK_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	thold_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCMRDPENDREQ_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMRDPENDREQ_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_PLBPPCMREARBITRATE_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMREARBITRATE_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMREQPRI_CPMPPCMPLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCMREQPRI_CPMPPCMPLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCMSSIZE_CPMPPCMPLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCMSSIZE_CPMPPCMPLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCMTIMEOUT_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMTIMEOUT_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMWRBTERM_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMWRBTERM_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMWRDACK_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMWRDACK_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCMWRPENDREQ_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCMWRPENDREQ_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0ABORT_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0ABORT_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	thold_PLBPPCS0BUSLOCK_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0BUSLOCK_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0LOCKERR_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0LOCKERR_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0MASTERID_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS0MASTERID_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS0MSIZE_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS0MSIZE_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS0PAVALID_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0PAVALID_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0RDBURST_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0RDBURST_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS0RDPENDREQ_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0RDPENDREQ_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0RDPRIM_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0RDPRIM_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0REQPRI_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS0REQPRI_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS0RNW_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0RNW_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0SAVALID_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0SAVALID_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0SIZE_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_PLBPPCS0SIZE_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	thold_PLBPPCS0TYPE_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 2) := (others => 0 ps);
	thold_PLBPPCS0TYPE_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 2) := (others => 0 ps);
	thold_PLBPPCS0UABUS_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(28 to 31) := (others => 0 ps);
	thold_PLBPPCS0UABUS_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(28 to 31) := (others => 0 ps);
	thold_PLBPPCS0WRBURST_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0WRBURST_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	thold_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS0WRPENDREQ_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0WRPENDREQ_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0WRPRIM_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS0WRPRIM_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1ABORT_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1ABORT_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	thold_PLBPPCS1BUSLOCK_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1BUSLOCK_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1LOCKERR_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1LOCKERR_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1MASTERID_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS1MASTERID_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS1MSIZE_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS1MSIZE_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS1PAVALID_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1PAVALID_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1RDBURST_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1RDBURST_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS1RDPENDREQ_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1RDPENDREQ_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1RDPRIM_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1RDPRIM_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1REQPRI_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS1REQPRI_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS1RNW_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1RNW_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1SAVALID_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1SAVALID_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1SIZE_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_PLBPPCS1SIZE_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	thold_PLBPPCS1TYPE_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 2) := (others => 0 ps);
	thold_PLBPPCS1TYPE_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 2) := (others => 0 ps);
	thold_PLBPPCS1UABUS_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(28 to 31) := (others => 0 ps);
	thold_PLBPPCS1UABUS_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(28 to 31) := (others => 0 ps);
	thold_PLBPPCS1WRBURST_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1WRBURST_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	thold_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	thold_PLBPPCS1WRPENDREQ_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1WRPENDREQ_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1WRPRIM_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_PLBPPCS1WRPRIM_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_TRCC440TRACEDISABLE_CPMC440CLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_TRCC440TRACEDISABLE_CPMC440CLK_posedge_posedge : VitalDelayType := 0 ps;
	thold_TRCC440TRIGGEREVENTIN_CPMC440CLK_negedge_posedge : VitalDelayType := 0 ps;
	thold_TRCC440TRIGGEREVENTIN_CPMC440CLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_CPMC440CORECLOCKINACTIVE_JTGC440TCK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_CPMC440CORECLOCKINACTIVE_JTGC440TCK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_CPMINTERCONNECTCLKNTO1_CPMINTERCONNECTCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_CPMINTERCONNECTCLKNTO1_CPMINTERCONNECTCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_DBGC440DEBUGHALT_CPMC440CLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_DBGC440DEBUGHALT_CPMC440CLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_DBGC440SYSTEMSTATUS_JTGC440TCK_negedge_posedge : VitalDelayArrayType(0 to 4) := (others => 0 ps);
	tsetup_DBGC440SYSTEMSTATUS_JTGC440TCK_posedge_posedge : VitalDelayArrayType(0 to 4) := (others => 0 ps);
	tsetup_DBGC440UNCONDDEBUGEVENT_CPMC440CLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_DBGC440UNCONDDEBUGEVENT_CPMC440CLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_DCRPPCDMACK_CPMDCRCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_DCRPPCDMACK_CPMDCRCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_DCRPPCDMTIMEOUTWAIT_CPMDCRCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_DCRPPCDMTIMEOUTWAIT_CPMDCRCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge : VitalDelayArrayType(0 to 9) := (others => 0 ps);
	tsetup_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge : VitalDelayArrayType(0 to 9) := (others => 0 ps);
	tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_DCRPPCDSREAD_CPMDCRCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_DCRPPCDSREAD_CPMDCRCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_DCRPPCDSWRITE_CPMDCRCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_DCRPPCDSWRITE_CPMDCRCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_FCMAPUCONFIRMINSTR_CPMFCMCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_FCMAPUCONFIRMINSTR_CPMFCMCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_FCMAPUCR_CPMFCMCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_FCMAPUCR_CPMFCMCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_FCMAPUDONE_CPMFCMCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_FCMAPUDONE_CPMFCMCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_FCMAPUEXCEPTION_CPMFCMCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_FCMAPUEXCEPTION_CPMFCMCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_FCMAPUFPSCRFEX_CPMFCMCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_FCMAPUFPSCRFEX_CPMFCMCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_FCMAPURESULTVALID_CPMFCMCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_FCMAPURESULTVALID_CPMFCMCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_FCMAPUSLEEPNOTREADY_CPMFCMCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_FCMAPUSLEEPNOTREADY_CPMFCMCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tsetup_JTGC440TDI_JTGC440TCK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_JTGC440TDI_JTGC440TCK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_JTGC440TMS_JTGC440TCK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_JTGC440TMS_JTGC440TCK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA0RSTENGINEREQ_CPMDMA0LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA0RSTENGINEREQ_CPMDMA0LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_LLDMA0RXEOFN_CPMDMA0LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA0RXEOFN_CPMDMA0LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA0RXEOPN_CPMDMA0LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA0RXEOPN_CPMDMA0LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA0RXREM_CPMDMA0LLCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_LLDMA0RXREM_CPMDMA0LLCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_LLDMA0RXSOFN_CPMDMA0LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA0RXSOFN_CPMDMA0LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA0RXSOPN_CPMDMA0LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA0RXSOPN_CPMDMA0LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA0RXSRCRDYN_CPMDMA0LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA0RXSRCRDYN_CPMDMA0LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA0TXDSTRDYN_CPMDMA0LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA0TXDSTRDYN_CPMDMA0LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA1RSTENGINEREQ_CPMDMA1LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA1RSTENGINEREQ_CPMDMA1LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_LLDMA1RXEOFN_CPMDMA1LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA1RXEOFN_CPMDMA1LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA1RXEOPN_CPMDMA1LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA1RXEOPN_CPMDMA1LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA1RXREM_CPMDMA1LLCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_LLDMA1RXREM_CPMDMA1LLCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_LLDMA1RXSOFN_CPMDMA1LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA1RXSOFN_CPMDMA1LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA1RXSOPN_CPMDMA1LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA1RXSOPN_CPMDMA1LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA1RXSRCRDYN_CPMDMA1LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA1RXSRCRDYN_CPMDMA1LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA1TXDSTRDYN_CPMDMA1LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA1TXDSTRDYN_CPMDMA1LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA2RSTENGINEREQ_CPMDMA2LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA2RSTENGINEREQ_CPMDMA2LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_LLDMA2RXEOFN_CPMDMA2LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA2RXEOFN_CPMDMA2LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA2RXEOPN_CPMDMA2LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA2RXEOPN_CPMDMA2LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA2RXREM_CPMDMA2LLCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_LLDMA2RXREM_CPMDMA2LLCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_LLDMA2RXSOFN_CPMDMA2LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA2RXSOFN_CPMDMA2LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA2RXSOPN_CPMDMA2LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA2RXSOPN_CPMDMA2LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA2RXSRCRDYN_CPMDMA2LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA2RXSRCRDYN_CPMDMA2LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA2TXDSTRDYN_CPMDMA2LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA2TXDSTRDYN_CPMDMA2LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA3RSTENGINEREQ_CPMDMA3LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA3RSTENGINEREQ_CPMDMA3LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_LLDMA3RXEOFN_CPMDMA3LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA3RXEOFN_CPMDMA3LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA3RXEOPN_CPMDMA3LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA3RXEOPN_CPMDMA3LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA3RXREM_CPMDMA3LLCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_LLDMA3RXREM_CPMDMA3LLCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_LLDMA3RXSOFN_CPMDMA3LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA3RXSOFN_CPMDMA3LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA3RXSOPN_CPMDMA3LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA3RXSOPN_CPMDMA3LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA3RXSRCRDYN_CPMDMA3LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA3RXSRCRDYN_CPMDMA3LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA3TXDSTRDYN_CPMDMA3LLCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_LLDMA3TXDSTRDYN_CPMDMA3LLCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_MCMIADDRREADYTOACCEPT_CPMMCCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_MCMIADDRREADYTOACCEPT_CPMMCCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_MCMIREADDATAERR_CPMMCCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_MCMIREADDATAERR_CPMMCCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_MCMIREADDATAVALID_CPMMCCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_MCMIREADDATAVALID_CPMMCCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tsetup_PLBPPCMADDRACK_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMADDRACK_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMMBUSY_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMMBUSY_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMMIRQ_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMMIRQ_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMMRDERR_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMMRDERR_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMMWRERR_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMMWRERR_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMRDBTERM_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMRDBTERM_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMRDDACK_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMRDDACK_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tsetup_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCMRDPENDREQ_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMRDPENDREQ_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_PLBPPCMREARBITRATE_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMREARBITRATE_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMREQPRI_CPMPPCMPLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCMREQPRI_CPMPPCMPLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCMSSIZE_CPMPPCMPLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCMSSIZE_CPMPPCMPLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCMTIMEOUT_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMTIMEOUT_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMWRBTERM_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMWRBTERM_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMWRDACK_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMWRDACK_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCMWRPENDREQ_CPMPPCMPLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCMWRPENDREQ_CPMPPCMPLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0ABORT_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0ABORT_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	tsetup_PLBPPCS0BUSLOCK_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0BUSLOCK_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0LOCKERR_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0LOCKERR_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0MASTERID_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS0MASTERID_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS0MSIZE_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS0MSIZE_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS0PAVALID_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0PAVALID_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0RDBURST_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0RDBURST_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS0RDPENDREQ_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0RDPENDREQ_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0RDPRIM_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0RDPRIM_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0REQPRI_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS0REQPRI_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS0RNW_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0RNW_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0SAVALID_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0SAVALID_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0SIZE_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_PLBPPCS0SIZE_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	tsetup_PLBPPCS0TYPE_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 2) := (others => 0 ps);
	tsetup_PLBPPCS0TYPE_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 2) := (others => 0 ps);
	tsetup_PLBPPCS0UABUS_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(28 to 31) := (others => 0 ps);
	tsetup_PLBPPCS0UABUS_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(28 to 31) := (others => 0 ps);
	tsetup_PLBPPCS0WRBURST_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0WRBURST_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tsetup_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS0WRPENDREQ_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0WRPENDREQ_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0WRPRIM_CPMPPCS0PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS0WRPRIM_CPMPPCS0PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1ABORT_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1ABORT_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	tsetup_PLBPPCS1BUSLOCK_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1BUSLOCK_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1LOCKERR_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1LOCKERR_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1MASTERID_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS1MASTERID_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS1MSIZE_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS1MSIZE_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS1PAVALID_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1PAVALID_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1RDBURST_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1RDBURST_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS1RDPENDREQ_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1RDPENDREQ_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1RDPRIM_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1RDPRIM_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1REQPRI_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS1REQPRI_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS1RNW_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1RNW_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1SAVALID_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1SAVALID_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1SIZE_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_PLBPPCS1SIZE_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	tsetup_PLBPPCS1TYPE_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 2) := (others => 0 ps);
	tsetup_PLBPPCS1TYPE_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 2) := (others => 0 ps);
	tsetup_PLBPPCS1UABUS_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(28 to 31) := (others => 0 ps);
	tsetup_PLBPPCS1UABUS_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(28 to 31) := (others => 0 ps);
	tsetup_PLBPPCS1WRBURST_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1WRBURST_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tsetup_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tsetup_PLBPPCS1WRPENDREQ_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1WRPENDREQ_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1WRPRIM_CPMPPCS1PLBCLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_PLBPPCS1WRPRIM_CPMPPCS1PLBCLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_TRCC440TRACEDISABLE_CPMC440CLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_TRCC440TRACEDISABLE_CPMC440CLK_posedge_posedge : VitalDelayType := 0 ps;
	tsetup_TRCC440TRIGGEREVENTIN_CPMC440CLK_negedge_posedge : VitalDelayType := 0 ps;
	tsetup_TRCC440TRIGGEREVENTIN_CPMC440CLK_posedge_posedge : VitalDelayType := 0 ps;

	ticd_CPMC440CLK : VitalDelayType := 0 ps;
	ticd_CPMDCRCLK : VitalDelayType := 0 ps;
	ticd_CPMDMA0LLCLK : VitalDelayType := 0 ps;
	ticd_CPMDMA1LLCLK : VitalDelayType := 0 ps;
	ticd_CPMDMA2LLCLK : VitalDelayType := 0 ps;
	ticd_CPMDMA3LLCLK : VitalDelayType := 0 ps;
	ticd_CPMFCMCLK : VitalDelayType := 0 ps;
	ticd_CPMINTERCONNECTCLK : VitalDelayType := 0 ps;
	ticd_CPMMCCLK : VitalDelayType := 0 ps;
	ticd_CPMPPCMPLBCLK : VitalDelayType := 0 ps;
	ticd_CPMPPCS0PLBCLK : VitalDelayType := 0 ps;
	ticd_CPMPPCS1PLBCLK : VitalDelayType := 0 ps;
	ticd_JTGC440TCK : VitalDelayType := 0 ps;

	tisd_CPMC440CORECLOCKINACTIVE_JTGC440TCK : VitalDelayType := 0 ps;
	tisd_CPMINTERCONNECTCLKNTO1_CPMINTERCONNECTCLK : VitalDelayType := 0 ps;
	tisd_DBGC440DEBUGHALT_CPMC440CLK : VitalDelayType := 0 ps;
	tisd_DBGC440SYSTEMSTATUS_JTGC440TCK : VitalDelayArrayType(0 to 4) := (others => 0 ps);
	tisd_DBGC440UNCONDDEBUGEVENT_CPMC440CLK : VitalDelayType := 0 ps;
	tisd_DCRPPCDMACK_CPMDCRCLK : VitalDelayType := 0 ps;
	tisd_DCRPPCDMDBUSIN_CPMDCRCLK : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tisd_DCRPPCDMTIMEOUTWAIT_CPMDCRCLK : VitalDelayType := 0 ps;
	tisd_DCRPPCDSABUS_CPMDCRCLK : VitalDelayArrayType(0 to 9) := (others => 0 ps);
	tisd_DCRPPCDSDBUSOUT_CPMDCRCLK : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tisd_DCRPPCDSREAD_CPMDCRCLK : VitalDelayType := 0 ps;
	tisd_DCRPPCDSWRITE_CPMDCRCLK : VitalDelayType := 0 ps;
	tisd_FCMAPUCONFIRMINSTR_CPMFCMCLK : VitalDelayType := 0 ps;
	tisd_FCMAPUCR_CPMFCMCLK : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tisd_FCMAPUDONE_CPMFCMCLK : VitalDelayType := 0 ps;
	tisd_FCMAPUEXCEPTION_CPMFCMCLK : VitalDelayType := 0 ps;
	tisd_FCMAPUFPSCRFEX_CPMFCMCLK : VitalDelayType := 0 ps;
	tisd_FCMAPURESULT_CPMFCMCLK : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tisd_FCMAPURESULTVALID_CPMFCMCLK : VitalDelayType := 0 ps;
	tisd_FCMAPUSLEEPNOTREADY_CPMFCMCLK : VitalDelayType := 0 ps;
	tisd_FCMAPUSTOREDATA_CPMFCMCLK : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tisd_JTGC440TDI_JTGC440TCK : VitalDelayType := 0 ps;
	tisd_JTGC440TMS_JTGC440TCK : VitalDelayType := 0 ps;
	tisd_LLDMA0RSTENGINEREQ_CPMDMA0LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA0RXD_CPMDMA0LLCLK : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tisd_LLDMA0RXEOFN_CPMDMA0LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA0RXEOPN_CPMDMA0LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA0RXREM_CPMDMA0LLCLK : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tisd_LLDMA0RXSOFN_CPMDMA0LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA0RXSOPN_CPMDMA0LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA0RXSRCRDYN_CPMDMA0LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA0TXDSTRDYN_CPMDMA0LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA1RSTENGINEREQ_CPMDMA1LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA1RXD_CPMDMA1LLCLK : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tisd_LLDMA1RXEOFN_CPMDMA1LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA1RXEOPN_CPMDMA1LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA1RXREM_CPMDMA1LLCLK : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tisd_LLDMA1RXSOFN_CPMDMA1LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA1RXSOPN_CPMDMA1LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA1RXSRCRDYN_CPMDMA1LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA1TXDSTRDYN_CPMDMA1LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA2RSTENGINEREQ_CPMDMA2LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA2RXD_CPMDMA2LLCLK : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tisd_LLDMA2RXEOFN_CPMDMA2LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA2RXEOPN_CPMDMA2LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA2RXREM_CPMDMA2LLCLK : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tisd_LLDMA2RXSOFN_CPMDMA2LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA2RXSOPN_CPMDMA2LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA2RXSRCRDYN_CPMDMA2LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA2TXDSTRDYN_CPMDMA2LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA3RSTENGINEREQ_CPMDMA3LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA3RXD_CPMDMA3LLCLK : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tisd_LLDMA3RXEOFN_CPMDMA3LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA3RXEOPN_CPMDMA3LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA3RXREM_CPMDMA3LLCLK : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tisd_LLDMA3RXSOFN_CPMDMA3LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA3RXSOPN_CPMDMA3LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA3RXSRCRDYN_CPMDMA3LLCLK : VitalDelayType := 0 ps;
	tisd_LLDMA3TXDSTRDYN_CPMDMA3LLCLK : VitalDelayType := 0 ps;
	tisd_MCMIADDRREADYTOACCEPT_CPMMCCLK : VitalDelayType := 0 ps;
	tisd_MCMIREADDATA_CPMMCCLK : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tisd_MCMIREADDATAERR_CPMMCCLK : VitalDelayType := 0 ps;
	tisd_MCMIREADDATAVALID_CPMMCCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCMADDRACK_CPMPPCMPLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCMMBUSY_CPMPPCMPLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCMMIRQ_CPMPPCMPLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCMMRDERR_CPMPPCMPLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCMMWRERR_CPMPPCMPLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCMRDBTERM_CPMPPCMPLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCMRDDACK_CPMPPCMPLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tisd_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tisd_PLBPPCMRDPENDREQ_CPMPPCMPLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCMRDWDADDR_CPMPPCMPLBCLK : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tisd_PLBPPCMREARBITRATE_CPMPPCMPLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCMREQPRI_CPMPPCMPLBCLK : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tisd_PLBPPCMSSIZE_CPMPPCMPLBCLK : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tisd_PLBPPCMTIMEOUT_CPMPPCMPLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCMWRBTERM_CPMPPCMPLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCMWRDACK_CPMPPCMPLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tisd_PLBPPCMWRPENDREQ_CPMPPCMPLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS0ABORT_CPMPPCS0PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tisd_PLBPPCS0BE_CPMPPCS0PLBCLK : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	tisd_PLBPPCS0BUSLOCK_CPMPPCS0PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS0LOCKERR_CPMPPCS0PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS0MASTERID_CPMPPCS0PLBCLK : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tisd_PLBPPCS0MSIZE_CPMPPCS0PLBCLK : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tisd_PLBPPCS0PAVALID_CPMPPCS0PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS0RDBURST_CPMPPCS0PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tisd_PLBPPCS0RDPENDREQ_CPMPPCS0PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS0RDPRIM_CPMPPCS0PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS0REQPRI_CPMPPCS0PLBCLK : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tisd_PLBPPCS0RNW_CPMPPCS0PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS0SAVALID_CPMPPCS0PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS0SIZE_CPMPPCS0PLBCLK : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	tisd_PLBPPCS0TYPE_CPMPPCS0PLBCLK : VitalDelayArrayType(0 to 2) := (others => 0 ps);
	tisd_PLBPPCS0UABUS_CPMPPCS0PLBCLK : VitalDelayArrayType(28 to 31) := (others => 0 ps);
	tisd_PLBPPCS0WRBURST_CPMPPCS0PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tisd_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tisd_PLBPPCS0WRPENDREQ_CPMPPCS0PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS0WRPRIM_CPMPPCS0PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS1ABORT_CPMPPCS1PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK : VitalDelayArrayType(0 to 31) := (others => 0 ps);
	tisd_PLBPPCS1BE_CPMPPCS1PLBCLK : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	tisd_PLBPPCS1BUSLOCK_CPMPPCS1PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS1LOCKERR_CPMPPCS1PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS1MASTERID_CPMPPCS1PLBCLK : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tisd_PLBPPCS1MSIZE_CPMPPCS1PLBCLK : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tisd_PLBPPCS1PAVALID_CPMPPCS1PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS1RDBURST_CPMPPCS1PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tisd_PLBPPCS1RDPENDREQ_CPMPPCS1PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS1RDPRIM_CPMPPCS1PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS1REQPRI_CPMPPCS1PLBCLK : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tisd_PLBPPCS1RNW_CPMPPCS1PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS1SAVALID_CPMPPCS1PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS1SIZE_CPMPPCS1PLBCLK : VitalDelayArrayType(0 to 3) := (others => 0 ps);
	tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK : VitalDelayArrayType(0 to 15) := (others => 0 ps);
	tisd_PLBPPCS1TYPE_CPMPPCS1PLBCLK : VitalDelayArrayType(0 to 2) := (others => 0 ps);
	tisd_PLBPPCS1UABUS_CPMPPCS1PLBCLK : VitalDelayArrayType(28 to 31) := (others => 0 ps);
	tisd_PLBPPCS1WRBURST_CPMPPCS1PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK : VitalDelayArrayType(0 to 127) := (others => 0 ps);
	tisd_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK : VitalDelayArrayType(0 to 1) := (others => 0 ps);
	tisd_PLBPPCS1WRPENDREQ_CPMPPCS1PLBCLK : VitalDelayType := 0 ps;
	tisd_PLBPPCS1WRPRIM_CPMPPCS1PLBCLK : VitalDelayType := 0 ps;
	tisd_TRCC440TRACEDISABLE_CPMC440CLK : VitalDelayType := 0 ps;
	tisd_TRCC440TRIGGEREVENTIN_CPMC440CLK : VitalDelayType := 0 ps 

  );

port (
		APUFCMDECFPUOP : out std_ulogic;
		APUFCMDECLDSTXFERSIZE : out std_logic_vector(0 to 2);
		APUFCMDECLOAD : out std_ulogic;
		APUFCMDECNONAUTON : out std_ulogic;
		APUFCMDECSTORE : out std_ulogic;
		APUFCMDECUDI : out std_logic_vector(0 to 3);
		APUFCMDECUDIVALID : out std_ulogic;
		APUFCMENDIAN : out std_ulogic;
		APUFCMFLUSH : out std_ulogic;
		APUFCMINSTRUCTION : out std_logic_vector(0 to 31);
		APUFCMINSTRVALID : out std_ulogic;
		APUFCMLOADBYTEADDR : out std_logic_vector(0 to 3);
		APUFCMLOADDATA : out std_logic_vector(0 to 127);
		APUFCMLOADDVALID : out std_ulogic;
		APUFCMMSRFE0 : out std_ulogic;
		APUFCMMSRFE1 : out std_ulogic;
		APUFCMNEXTINSTRREADY : out std_ulogic;
		APUFCMOPERANDVALID : out std_ulogic;
		APUFCMRADATA : out std_logic_vector(0 to 31);
		APUFCMRBDATA : out std_logic_vector(0 to 31);
		APUFCMWRITEBACKOK : out std_ulogic;
		C440CPMCORESLEEPREQ : out std_ulogic;
		C440CPMDECIRPTREQ : out std_ulogic;
		C440CPMFITIRPTREQ : out std_ulogic;
		C440CPMMSRCE : out std_ulogic;
		C440CPMMSREE : out std_ulogic;
		C440CPMTIMERRESETREQ : out std_ulogic;
		C440CPMWDIRPTREQ : out std_ulogic;
		C440DBGSYSTEMCONTROL : out std_logic_vector(0 to 7);
		C440JTGTDO : out std_ulogic;
		C440JTGTDOEN : out std_ulogic;
		C440MACHINECHECK : out std_ulogic;
		C440RSTCHIPRESETREQ : out std_ulogic;
		C440RSTCORERESETREQ : out std_ulogic;
		C440RSTSYSTEMRESETREQ : out std_ulogic;
		C440TRCBRANCHSTATUS : out std_logic_vector(0 to 2);
		C440TRCCYCLE : out std_ulogic;
		C440TRCEXECUTIONSTATUS : out std_logic_vector(0 to 4);
		C440TRCTRACESTATUS : out std_logic_vector(0 to 6);
		C440TRCTRIGGEREVENTOUT : out std_ulogic;
		C440TRCTRIGGEREVENTTYPE : out std_logic_vector(0 to 13);
		DMA0LLRSTENGINEACK : out std_ulogic;
		DMA0LLRXDSTRDYN : out std_ulogic;
		DMA0LLTXD : out std_logic_vector(0 to 31);
		DMA0LLTXEOFN : out std_ulogic;
		DMA0LLTXEOPN : out std_ulogic;
		DMA0LLTXREM : out std_logic_vector(0 to 3);
		DMA0LLTXSOFN : out std_ulogic;
		DMA0LLTXSOPN : out std_ulogic;
		DMA0LLTXSRCRDYN : out std_ulogic;
		DMA0RXIRQ : out std_ulogic;
		DMA0TXIRQ : out std_ulogic;
		DMA1LLRSTENGINEACK : out std_ulogic;
		DMA1LLRXDSTRDYN : out std_ulogic;
		DMA1LLTXD : out std_logic_vector(0 to 31);
		DMA1LLTXEOFN : out std_ulogic;
		DMA1LLTXEOPN : out std_ulogic;
		DMA1LLTXREM : out std_logic_vector(0 to 3);
		DMA1LLTXSOFN : out std_ulogic;
		DMA1LLTXSOPN : out std_ulogic;
		DMA1LLTXSRCRDYN : out std_ulogic;
		DMA1RXIRQ : out std_ulogic;
		DMA1TXIRQ : out std_ulogic;
		DMA2LLRSTENGINEACK : out std_ulogic;
		DMA2LLRXDSTRDYN : out std_ulogic;
		DMA2LLTXD : out std_logic_vector(0 to 31);
		DMA2LLTXEOFN : out std_ulogic;
		DMA2LLTXEOPN : out std_ulogic;
		DMA2LLTXREM : out std_logic_vector(0 to 3);
		DMA2LLTXSOFN : out std_ulogic;
		DMA2LLTXSOPN : out std_ulogic;
		DMA2LLTXSRCRDYN : out std_ulogic;
		DMA2RXIRQ : out std_ulogic;
		DMA2TXIRQ : out std_ulogic;
		DMA3LLRSTENGINEACK : out std_ulogic;
		DMA3LLRXDSTRDYN : out std_ulogic;
		DMA3LLTXD : out std_logic_vector(0 to 31);
		DMA3LLTXEOFN : out std_ulogic;
		DMA3LLTXEOPN : out std_ulogic;
		DMA3LLTXREM : out std_logic_vector(0 to 3);
		DMA3LLTXSOFN : out std_ulogic;
		DMA3LLTXSOPN : out std_ulogic;
		DMA3LLTXSRCRDYN : out std_ulogic;
		DMA3RXIRQ : out std_ulogic;
		DMA3TXIRQ : out std_ulogic;
		MIMCADDRESS : out std_logic_vector(0 to 35);
		MIMCADDRESSVALID : out std_ulogic;
		MIMCBANKCONFLICT : out std_ulogic;
		MIMCBYTEENABLE : out std_logic_vector(0 to 15);
		MIMCREADNOTWRITE : out std_ulogic;
		MIMCROWCONFLICT : out std_ulogic;
		MIMCWRITEDATA : out std_logic_vector(0 to 127);
		MIMCWRITEDATAVALID : out std_ulogic;
		PPCCPMINTERCONNECTBUSY : out std_ulogic;
		PPCDMDCRABUS : out std_logic_vector(0 to 9);
		PPCDMDCRDBUSOUT : out std_logic_vector(0 to 31);
		PPCDMDCRREAD : out std_ulogic;
		PPCDMDCRUABUS : out std_logic_vector(20 to 21);
		PPCDMDCRWRITE : out std_ulogic;
		PPCDSDCRACK : out std_ulogic;
		PPCDSDCRDBUSIN : out std_logic_vector(0 to 31);
		PPCDSDCRTIMEOUTWAIT : out std_ulogic;
		PPCEICINTERCONNECTIRQ : out std_ulogic;
		PPCMPLBABORT : out std_ulogic;
		PPCMPLBABUS : out std_logic_vector(0 to 31);
		PPCMPLBBE : out std_logic_vector(0 to 15);
		PPCMPLBBUSLOCK : out std_ulogic;
		PPCMPLBLOCKERR : out std_ulogic;
		PPCMPLBPRIORITY : out std_logic_vector(0 to 1);
		PPCMPLBRDBURST : out std_ulogic;
		PPCMPLBREQUEST : out std_ulogic;
		PPCMPLBRNW : out std_ulogic;
		PPCMPLBSIZE : out std_logic_vector(0 to 3);
		PPCMPLBTATTRIBUTE : out std_logic_vector(0 to 15);
		PPCMPLBTYPE : out std_logic_vector(0 to 2);
		PPCMPLBUABUS : out std_logic_vector(28 to 31);
		PPCMPLBWRBURST : out std_ulogic;
		PPCMPLBWRDBUS : out std_logic_vector(0 to 127);
		PPCS0PLBADDRACK : out std_ulogic;
		PPCS0PLBMBUSY : out std_logic_vector(0 to 3);
		PPCS0PLBMIRQ : out std_logic_vector(0 to 3);
		PPCS0PLBMRDERR : out std_logic_vector(0 to 3);
		PPCS0PLBMWRERR : out std_logic_vector(0 to 3);
		PPCS0PLBRDBTERM : out std_ulogic;
		PPCS0PLBRDCOMP : out std_ulogic;
		PPCS0PLBRDDACK : out std_ulogic;
		PPCS0PLBRDDBUS : out std_logic_vector(0 to 127);
		PPCS0PLBRDWDADDR : out std_logic_vector(0 to 3);
		PPCS0PLBREARBITRATE : out std_ulogic;
		PPCS0PLBSSIZE : out std_logic_vector(0 to 1);
		PPCS0PLBWAIT : out std_ulogic;
		PPCS0PLBWRBTERM : out std_ulogic;
		PPCS0PLBWRCOMP : out std_ulogic;
		PPCS0PLBWRDACK : out std_ulogic;
		PPCS1PLBADDRACK : out std_ulogic;
		PPCS1PLBMBUSY : out std_logic_vector(0 to 3);
		PPCS1PLBMIRQ : out std_logic_vector(0 to 3);
		PPCS1PLBMRDERR : out std_logic_vector(0 to 3);
		PPCS1PLBMWRERR : out std_logic_vector(0 to 3);
		PPCS1PLBRDBTERM : out std_ulogic;
		PPCS1PLBRDCOMP : out std_ulogic;
		PPCS1PLBRDDACK : out std_ulogic;
		PPCS1PLBRDDBUS : out std_logic_vector(0 to 127);
		PPCS1PLBRDWDADDR : out std_logic_vector(0 to 3);
		PPCS1PLBREARBITRATE : out std_ulogic;
		PPCS1PLBSSIZE : out std_logic_vector(0 to 1);
		PPCS1PLBWAIT : out std_ulogic;
		PPCS1PLBWRBTERM : out std_ulogic;
		PPCS1PLBWRCOMP : out std_ulogic;
		PPCS1PLBWRDACK : out std_ulogic;

		CPMC440CLK : in std_ulogic;
		CPMC440CLKEN : in std_ulogic;
		CPMC440CORECLOCKINACTIVE : in std_ulogic;
		CPMC440TIMERCLOCK : in std_ulogic;
		CPMDCRCLK : in std_ulogic;
		CPMDMA0LLCLK : in std_ulogic;
		CPMDMA1LLCLK : in std_ulogic;
		CPMDMA2LLCLK : in std_ulogic;
		CPMDMA3LLCLK : in std_ulogic;
		CPMFCMCLK : in std_ulogic;
		CPMINTERCONNECTCLK : in std_ulogic;
		CPMINTERCONNECTCLKEN : in std_ulogic;
		CPMINTERCONNECTCLKNTO1 : in std_ulogic;
		CPMMCCLK : in std_ulogic;
		CPMPPCMPLBCLK : in std_ulogic;
		CPMPPCS0PLBCLK : in std_ulogic;
		CPMPPCS1PLBCLK : in std_ulogic;
		DBGC440DEBUGHALT : in std_ulogic;
		DBGC440SYSTEMSTATUS : in std_logic_vector(0 to 4);
		DBGC440UNCONDDEBUGEVENT : in std_ulogic;
		DCRPPCDMACK : in std_ulogic;
		DCRPPCDMDBUSIN : in std_logic_vector(0 to 31);
		DCRPPCDMTIMEOUTWAIT : in std_ulogic;
		DCRPPCDSABUS : in std_logic_vector(0 to 9);
		DCRPPCDSDBUSOUT : in std_logic_vector(0 to 31);
		DCRPPCDSREAD : in std_ulogic;
		DCRPPCDSWRITE : in std_ulogic;
		EICC440CRITIRQ : in std_ulogic;
		EICC440EXTIRQ : in std_ulogic;
		FCMAPUCONFIRMINSTR : in std_ulogic;
		FCMAPUCR : in std_logic_vector(0 to 3);
		FCMAPUDONE : in std_ulogic;
		FCMAPUEXCEPTION : in std_ulogic;
		FCMAPUFPSCRFEX : in std_ulogic;
		FCMAPURESULT : in std_logic_vector(0 to 31);
		FCMAPURESULTVALID : in std_ulogic;
		FCMAPUSLEEPNOTREADY : in std_ulogic;
		FCMAPUSTOREDATA : in std_logic_vector(0 to 127);
		JTGC440TCK : in std_ulogic;
		JTGC440TDI : in std_ulogic;
		JTGC440TMS : in std_ulogic;
		JTGC440TRSTNEG : in std_ulogic;
		LLDMA0RSTENGINEREQ : in std_ulogic;
		LLDMA0RXD : in std_logic_vector(0 to 31);
		LLDMA0RXEOFN : in std_ulogic;
		LLDMA0RXEOPN : in std_ulogic;
		LLDMA0RXREM : in std_logic_vector(0 to 3);
		LLDMA0RXSOFN : in std_ulogic;
		LLDMA0RXSOPN : in std_ulogic;
		LLDMA0RXSRCRDYN : in std_ulogic;
		LLDMA0TXDSTRDYN : in std_ulogic;
		LLDMA1RSTENGINEREQ : in std_ulogic;
		LLDMA1RXD : in std_logic_vector(0 to 31);
		LLDMA1RXEOFN : in std_ulogic;
		LLDMA1RXEOPN : in std_ulogic;
		LLDMA1RXREM : in std_logic_vector(0 to 3);
		LLDMA1RXSOFN : in std_ulogic;
		LLDMA1RXSOPN : in std_ulogic;
		LLDMA1RXSRCRDYN : in std_ulogic;
		LLDMA1TXDSTRDYN : in std_ulogic;
		LLDMA2RSTENGINEREQ : in std_ulogic;
		LLDMA2RXD : in std_logic_vector(0 to 31);
		LLDMA2RXEOFN : in std_ulogic;
		LLDMA2RXEOPN : in std_ulogic;
		LLDMA2RXREM : in std_logic_vector(0 to 3);
		LLDMA2RXSOFN : in std_ulogic;
		LLDMA2RXSOPN : in std_ulogic;
		LLDMA2RXSRCRDYN : in std_ulogic;
		LLDMA2TXDSTRDYN : in std_ulogic;
		LLDMA3RSTENGINEREQ : in std_ulogic;
		LLDMA3RXD : in std_logic_vector(0 to 31);
		LLDMA3RXEOFN : in std_ulogic;
		LLDMA3RXEOPN : in std_ulogic;
		LLDMA3RXREM : in std_logic_vector(0 to 3);
		LLDMA3RXSOFN : in std_ulogic;
		LLDMA3RXSOPN : in std_ulogic;
		LLDMA3RXSRCRDYN : in std_ulogic;
		LLDMA3TXDSTRDYN : in std_ulogic;
		MCMIADDRREADYTOACCEPT : in std_ulogic;
		MCMIREADDATA : in std_logic_vector(0 to 127);
		MCMIREADDATAERR : in std_ulogic;
		MCMIREADDATAVALID : in std_ulogic;
		PLBPPCMADDRACK : in std_ulogic;
		PLBPPCMMBUSY : in std_ulogic;
		PLBPPCMMIRQ : in std_ulogic;
		PLBPPCMMRDERR : in std_ulogic;
		PLBPPCMMWRERR : in std_ulogic;
		PLBPPCMRDBTERM : in std_ulogic;
		PLBPPCMRDDACK : in std_ulogic;
		PLBPPCMRDDBUS : in std_logic_vector(0 to 127);
		PLBPPCMRDPENDPRI : in std_logic_vector(0 to 1);
		PLBPPCMRDPENDREQ : in std_ulogic;
		PLBPPCMRDWDADDR : in std_logic_vector(0 to 3);
		PLBPPCMREARBITRATE : in std_ulogic;
		PLBPPCMREQPRI : in std_logic_vector(0 to 1);
		PLBPPCMSSIZE : in std_logic_vector(0 to 1);
		PLBPPCMTIMEOUT : in std_ulogic;
		PLBPPCMWRBTERM : in std_ulogic;
		PLBPPCMWRDACK : in std_ulogic;
		PLBPPCMWRPENDPRI : in std_logic_vector(0 to 1);
		PLBPPCMWRPENDREQ : in std_ulogic;
		PLBPPCS0ABORT : in std_ulogic;
		PLBPPCS0ABUS : in std_logic_vector(0 to 31);
		PLBPPCS0BE : in std_logic_vector(0 to 15);
		PLBPPCS0BUSLOCK : in std_ulogic;
		PLBPPCS0LOCKERR : in std_ulogic;
		PLBPPCS0MASTERID : in std_logic_vector(0 to 1);
		PLBPPCS0MSIZE : in std_logic_vector(0 to 1);
		PLBPPCS0PAVALID : in std_ulogic;
		PLBPPCS0RDBURST : in std_ulogic;
		PLBPPCS0RDPENDPRI : in std_logic_vector(0 to 1);
		PLBPPCS0RDPENDREQ : in std_ulogic;
		PLBPPCS0RDPRIM : in std_ulogic;
		PLBPPCS0REQPRI : in std_logic_vector(0 to 1);
		PLBPPCS0RNW : in std_ulogic;
		PLBPPCS0SAVALID : in std_ulogic;
		PLBPPCS0SIZE : in std_logic_vector(0 to 3);
		PLBPPCS0TATTRIBUTE : in std_logic_vector(0 to 15);
		PLBPPCS0TYPE : in std_logic_vector(0 to 2);
		PLBPPCS0UABUS : in std_logic_vector(28 to 31);
		PLBPPCS0WRBURST : in std_ulogic;
		PLBPPCS0WRDBUS : in std_logic_vector(0 to 127);
		PLBPPCS0WRPENDPRI : in std_logic_vector(0 to 1);
		PLBPPCS0WRPENDREQ : in std_ulogic;
		PLBPPCS0WRPRIM : in std_ulogic;
		PLBPPCS1ABORT : in std_ulogic;
		PLBPPCS1ABUS : in std_logic_vector(0 to 31);
		PLBPPCS1BE : in std_logic_vector(0 to 15);
		PLBPPCS1BUSLOCK : in std_ulogic;
		PLBPPCS1LOCKERR : in std_ulogic;
		PLBPPCS1MASTERID : in std_logic_vector(0 to 1);
		PLBPPCS1MSIZE : in std_logic_vector(0 to 1);
		PLBPPCS1PAVALID : in std_ulogic;
		PLBPPCS1RDBURST : in std_ulogic;
		PLBPPCS1RDPENDPRI : in std_logic_vector(0 to 1);
		PLBPPCS1RDPENDREQ : in std_ulogic;
		PLBPPCS1RDPRIM : in std_ulogic;
		PLBPPCS1REQPRI : in std_logic_vector(0 to 1);
		PLBPPCS1RNW : in std_ulogic;
		PLBPPCS1SAVALID : in std_ulogic;
		PLBPPCS1SIZE : in std_logic_vector(0 to 3);
		PLBPPCS1TATTRIBUTE : in std_logic_vector(0 to 15);
		PLBPPCS1TYPE : in std_logic_vector(0 to 2);
		PLBPPCS1UABUS : in std_logic_vector(28 to 31);
		PLBPPCS1WRBURST : in std_ulogic;
		PLBPPCS1WRDBUS : in std_logic_vector(0 to 127);
		PLBPPCS1WRPENDPRI : in std_logic_vector(0 to 1);
		PLBPPCS1WRPENDREQ : in std_ulogic;
		PLBPPCS1WRPRIM : in std_ulogic;
		RSTC440RESETCHIP : in std_ulogic;
		RSTC440RESETCORE : in std_ulogic;
		RSTC440RESETSYSTEM : in std_ulogic;
		TIEC440DCURDLDCACHEPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440DCURDNONCACHEPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440DCURDTOUCHPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440DCURDURGENTPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440DCUWRFLUSHPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440DCUWRSTOREPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440DCUWRURGENTPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440ENDIANRESET : in std_ulogic;
		TIEC440ERPNRESET : in std_logic_vector(0 to 3);
		TIEC440ICURDFETCHPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440ICURDSPECPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440ICURDTOUCHPLBPRIO : in std_logic_vector(0 to 1);
		TIEC440PIR : in std_logic_vector(28 to 31);
		TIEC440PVR : in std_logic_vector(28 to 31);
		TIEC440USERRESET : in std_logic_vector(0 to 3);
		TIEDCRBASEADDR : in std_logic_vector(0 to 1);
		TRCC440TRACEDISABLE : in std_ulogic;
		TRCC440TRIGGEREVENTIN : in std_ulogic
     );
attribute VITAL_LEVEL0 of X_PPC440 :     entity is true;

end X_PPC440;

architecture X_PPC440_V of X_PPC440 is

  component PPC440_SWIFT
    port (
      APUFCMDECFPUOP       : out std_ulogic;
      APUFCMDECLDSTXFERSIZE : out std_logic_vector(0 to 2);
      APUFCMDECLOAD        : out std_ulogic;
      APUFCMDECNONAUTON    : out std_ulogic;
      APUFCMDECSTORE       : out std_ulogic;
      APUFCMDECUDI         : out std_logic_vector(0 to 3);
      APUFCMDECUDIVALID    : out std_ulogic;
      APUFCMENDIAN         : out std_ulogic;
      APUFCMFLUSH          : out std_ulogic;
      APUFCMINSTRUCTION    : out std_logic_vector(0 to 31);
      APUFCMINSTRVALID     : out std_ulogic;
      APUFCMLOADBYTEADDR   : out std_logic_vector(0 to 3);
      APUFCMLOADDATA       : out std_logic_vector(0 to 127);
      APUFCMLOADDVALID     : out std_ulogic;
      APUFCMMSRFE0         : out std_ulogic;
      APUFCMMSRFE1         : out std_ulogic;
      APUFCMNEXTINSTRREADY : out std_ulogic;
      APUFCMOPERANDVALID   : out std_ulogic;
      APUFCMRADATA         : out std_logic_vector(0 to 31);
      APUFCMRBDATA         : out std_logic_vector(0 to 31);
      APUFCMWRITEBACKOK    : out std_ulogic;
      C440CPMCORESLEEPREQ  : out std_ulogic;
      C440CPMDECIRPTREQ    : out std_ulogic;
      C440CPMFITIRPTREQ    : out std_ulogic;
      C440CPMMSRCE         : out std_ulogic;
      C440CPMMSREE         : out std_ulogic;
      C440CPMTIMERRESETREQ : out std_ulogic;
      C440CPMWDIRPTREQ     : out std_ulogic;
      C440DBGSYSTEMCONTROL : out std_logic_vector(0 to 7);
      C440JTGTDO           : out std_ulogic;
      C440JTGTDOEN         : out std_ulogic;
      C440MACHINECHECK     : out std_ulogic;
      C440RSTCHIPRESETREQ  : out std_ulogic;
      C440RSTCORERESETREQ  : out std_ulogic;
      C440RSTSYSTEMRESETREQ : out std_ulogic;
      C440TRCBRANCHSTATUS  : out std_logic_vector(0 to 2);
      C440TRCCYCLE         : out std_ulogic;
      C440TRCEXECUTIONSTATUS : out std_logic_vector(0 to 4);
      C440TRCTRACESTATUS   : out std_logic_vector(0 to 6);
      C440TRCTRIGGEREVENTOUT : out std_ulogic;
      C440TRCTRIGGEREVENTTYPE : out std_logic_vector(0 to 13);
      DMA0LLRSTENGINEACK   : out std_ulogic;
      DMA0LLRXDSTRDYN      : out std_ulogic;
      DMA0LLTXD            : out std_logic_vector(0 to 31);
      DMA0LLTXEOFN         : out std_ulogic;
      DMA0LLTXEOPN         : out std_ulogic;
      DMA0LLTXREM          : out std_logic_vector(0 to 3);
      DMA0LLTXSOFN         : out std_ulogic;
      DMA0LLTXSOPN         : out std_ulogic;
      DMA0LLTXSRCRDYN      : out std_ulogic;
      DMA0RXIRQ            : out std_ulogic;
      DMA0TXIRQ            : out std_ulogic;
      DMA1LLRSTENGINEACK   : out std_ulogic;
      DMA1LLRXDSTRDYN      : out std_ulogic;
      DMA1LLTXD            : out std_logic_vector(0 to 31);
      DMA1LLTXEOFN         : out std_ulogic;
      DMA1LLTXEOPN         : out std_ulogic;
      DMA1LLTXREM          : out std_logic_vector(0 to 3);
      DMA1LLTXSOFN         : out std_ulogic;
      DMA1LLTXSOPN         : out std_ulogic;
      DMA1LLTXSRCRDYN      : out std_ulogic;
      DMA1RXIRQ            : out std_ulogic;
      DMA1TXIRQ            : out std_ulogic;
      DMA2LLRSTENGINEACK   : out std_ulogic;
      DMA2LLRXDSTRDYN      : out std_ulogic;
      DMA2LLTXD            : out std_logic_vector(0 to 31);
      DMA2LLTXEOFN         : out std_ulogic;
      DMA2LLTXEOPN         : out std_ulogic;
      DMA2LLTXREM          : out std_logic_vector(0 to 3);
      DMA2LLTXSOFN         : out std_ulogic;
      DMA2LLTXSOPN         : out std_ulogic;
      DMA2LLTXSRCRDYN      : out std_ulogic;
      DMA2RXIRQ            : out std_ulogic;
      DMA2TXIRQ            : out std_ulogic;
      DMA3LLRSTENGINEACK   : out std_ulogic;
      DMA3LLRXDSTRDYN      : out std_ulogic;
      DMA3LLTXD            : out std_logic_vector(0 to 31);
      DMA3LLTXEOFN         : out std_ulogic;
      DMA3LLTXEOPN         : out std_ulogic;
      DMA3LLTXREM          : out std_logic_vector(0 to 3);
      DMA3LLTXSOFN         : out std_ulogic;
      DMA3LLTXSOPN         : out std_ulogic;
      DMA3LLTXSRCRDYN      : out std_ulogic;
      DMA3RXIRQ            : out std_ulogic;
      DMA3TXIRQ            : out std_ulogic;
      MIMCADDRESS          : out std_logic_vector(0 to 35);
      MIMCADDRESSVALID     : out std_ulogic;
      MIMCBANKCONFLICT     : out std_ulogic;
      MIMCBYTEENABLE       : out std_logic_vector(0 to 15);
      MIMCREADNOTWRITE     : out std_ulogic;
      MIMCROWCONFLICT      : out std_ulogic;
      MIMCWRITEDATA        : out std_logic_vector(0 to 127);
      MIMCWRITEDATAVALID   : out std_ulogic;
      PPCCPMINTERCONNECTBUSY : out std_ulogic;
      PPCDMDCRABUS         : out std_logic_vector(0 to 9);
      PPCDMDCRDBUSOUT      : out std_logic_vector(0 to 31);
      PPCDMDCRREAD         : out std_ulogic;
      PPCDMDCRUABUS        : out std_logic_vector(20 to 21);
      PPCDMDCRWRITE        : out std_ulogic;
      PPCDSDCRACK          : out std_ulogic;
      PPCDSDCRDBUSIN       : out std_logic_vector(0 to 31);
      PPCDSDCRTIMEOUTWAIT  : out std_ulogic;
      PPCEICINTERCONNECTIRQ : out std_ulogic;
      PPCMPLBABORT         : out std_ulogic;
      PPCMPLBABUS          : out std_logic_vector(0 to 31);
      PPCMPLBBE            : out std_logic_vector(0 to 15);
      PPCMPLBBUSLOCK       : out std_ulogic;
      PPCMPLBLOCKERR       : out std_ulogic;
      PPCMPLBPRIORITY      : out std_logic_vector(0 to 1);
      PPCMPLBRDBURST       : out std_ulogic;
      PPCMPLBREQUEST       : out std_ulogic;
      PPCMPLBRNW           : out std_ulogic;
      PPCMPLBSIZE          : out std_logic_vector(0 to 3);
      PPCMPLBTATTRIBUTE    : out std_logic_vector(0 to 15);
      PPCMPLBTYPE          : out std_logic_vector(0 to 2);
      PPCMPLBUABUS         : out std_logic_vector(28 to 31);
      PPCMPLBWRBURST       : out std_ulogic;
      PPCMPLBWRDBUS        : out std_logic_vector(0 to 127);
      PPCS0PLBADDRACK      : out std_ulogic;
      PPCS0PLBMBUSY        : out std_logic_vector(0 to 3);
      PPCS0PLBMIRQ         : out std_logic_vector(0 to 3);
      PPCS0PLBMRDERR       : out std_logic_vector(0 to 3);
      PPCS0PLBMWRERR       : out std_logic_vector(0 to 3);
      PPCS0PLBRDBTERM      : out std_ulogic;
      PPCS0PLBRDCOMP       : out std_ulogic;
      PPCS0PLBRDDACK       : out std_ulogic;
      PPCS0PLBRDDBUS       : out std_logic_vector(0 to 127);
      PPCS0PLBRDWDADDR     : out std_logic_vector(0 to 3);
      PPCS0PLBREARBITRATE  : out std_ulogic;
      PPCS0PLBSSIZE        : out std_logic_vector(0 to 1);
      PPCS0PLBWAIT         : out std_ulogic;
      PPCS0PLBWRBTERM      : out std_ulogic;
      PPCS0PLBWRCOMP       : out std_ulogic;
      PPCS0PLBWRDACK       : out std_ulogic;
      PPCS1PLBADDRACK      : out std_ulogic;
      PPCS1PLBMBUSY        : out std_logic_vector(0 to 3);
      PPCS1PLBMIRQ         : out std_logic_vector(0 to 3);
      PPCS1PLBMRDERR       : out std_logic_vector(0 to 3);
      PPCS1PLBMWRERR       : out std_logic_vector(0 to 3);
      PPCS1PLBRDBTERM      : out std_ulogic;
      PPCS1PLBRDCOMP       : out std_ulogic;
      PPCS1PLBRDDACK       : out std_ulogic;
      PPCS1PLBRDDBUS       : out std_logic_vector(0 to 127);
      PPCS1PLBRDWDADDR     : out std_logic_vector(0 to 3);
      PPCS1PLBREARBITRATE  : out std_ulogic;
      PPCS1PLBSSIZE        : out std_logic_vector(0 to 1);
      PPCS1PLBWAIT         : out std_ulogic;
      PPCS1PLBWRBTERM      : out std_ulogic;
      PPCS1PLBWRCOMP       : out std_ulogic;
      PPCS1PLBWRDACK       : out std_ulogic;

      CPMC440CLK           : in std_ulogic;
      CPMC440CLKEN         : in std_ulogic;
      CPMC440CORECLOCKINACTIVE : in std_ulogic;
      CPMC440TIMERCLOCK    : in std_ulogic;
      CPMDCRCLK            : in std_ulogic;
      CPMDMA0LLCLK         : in std_ulogic;
      CPMDMA1LLCLK         : in std_ulogic;
      CPMDMA2LLCLK         : in std_ulogic;
      CPMDMA3LLCLK         : in std_ulogic;
      CPMFCMCLK            : in std_ulogic;
      CPMINTERCONNECTCLK   : in std_ulogic;
      CPMINTERCONNECTCLKEN : in std_ulogic;
      CPMINTERCONNECTCLKNTO1 : in std_ulogic;
      CPMMCCLK             : in std_ulogic;
      CPMPPCMPLBCLK        : in std_ulogic;
      CPMPPCS0PLBCLK       : in std_ulogic;
      CPMPPCS1PLBCLK       : in std_ulogic;
      DBGC440DEBUGHALT     : in std_ulogic;
      DBGC440SYSTEMSTATUS  : in std_logic_vector(0 to 4);
      DBGC440UNCONDDEBUGEVENT : in std_ulogic;
      DCRPPCDMACK          : in std_ulogic;
      DCRPPCDMDBUSIN       : in std_logic_vector(0 to 31);
      DCRPPCDMTIMEOUTWAIT  : in std_ulogic;
      DCRPPCDSABUS         : in std_logic_vector(0 to 9);
      DCRPPCDSDBUSOUT      : in std_logic_vector(0 to 31);
      DCRPPCDSREAD         : in std_ulogic;
      DCRPPCDSWRITE        : in std_ulogic;
      EICC440CRITIRQ       : in std_ulogic;
      EICC440EXTIRQ        : in std_ulogic;
      FCMAPUCONFIRMINSTR   : in std_ulogic;
      FCMAPUCR             : in std_logic_vector(0 to 3);
      FCMAPUDONE           : in std_ulogic;
      FCMAPUEXCEPTION      : in std_ulogic;
      FCMAPUFPSCRFEX       : in std_ulogic;
      FCMAPURESULT         : in std_logic_vector(0 to 31);
      FCMAPURESULTVALID    : in std_ulogic;
      FCMAPUSLEEPNOTREADY  : in std_ulogic;
      FCMAPUSTOREDATA      : in std_logic_vector(0 to 127);
      GSR                  : in std_ulogic;
      JTGC440TCK           : in std_ulogic;
      JTGC440TDI           : in std_ulogic;
      JTGC440TMS           : in std_ulogic;
      JTGC440TRSTNEG       : in std_ulogic;
      LLDMA0RSTENGINEREQ   : in std_ulogic;
      LLDMA0RXD            : in std_logic_vector(0 to 31);
      LLDMA0RXEOFN         : in std_ulogic;
      LLDMA0RXEOPN         : in std_ulogic;
      LLDMA0RXREM          : in std_logic_vector(0 to 3);
      LLDMA0RXSOFN         : in std_ulogic;
      LLDMA0RXSOPN         : in std_ulogic;
      LLDMA0RXSRCRDYN      : in std_ulogic;
      LLDMA0TXDSTRDYN      : in std_ulogic;
      LLDMA1RSTENGINEREQ   : in std_ulogic;
      LLDMA1RXD            : in std_logic_vector(0 to 31);
      LLDMA1RXEOFN         : in std_ulogic;
      LLDMA1RXEOPN         : in std_ulogic;
      LLDMA1RXREM          : in std_logic_vector(0 to 3);
      LLDMA1RXSOFN         : in std_ulogic;
      LLDMA1RXSOPN         : in std_ulogic;
      LLDMA1RXSRCRDYN      : in std_ulogic;
      LLDMA1TXDSTRDYN      : in std_ulogic;
      LLDMA2RSTENGINEREQ   : in std_ulogic;
      LLDMA2RXD            : in std_logic_vector(0 to 31);
      LLDMA2RXEOFN         : in std_ulogic;
      LLDMA2RXEOPN         : in std_ulogic;
      LLDMA2RXREM          : in std_logic_vector(0 to 3);
      LLDMA2RXSOFN         : in std_ulogic;
      LLDMA2RXSOPN         : in std_ulogic;
      LLDMA2RXSRCRDYN      : in std_ulogic;
      LLDMA2TXDSTRDYN      : in std_ulogic;
      LLDMA3RSTENGINEREQ   : in std_ulogic;
      LLDMA3RXD            : in std_logic_vector(0 to 31);
      LLDMA3RXEOFN         : in std_ulogic;
      LLDMA3RXEOPN         : in std_ulogic;
      LLDMA3RXREM          : in std_logic_vector(0 to 3);
      LLDMA3RXSOFN         : in std_ulogic;
      LLDMA3RXSOPN         : in std_ulogic;
      LLDMA3RXSRCRDYN      : in std_ulogic;
      LLDMA3TXDSTRDYN      : in std_ulogic;
      MCMIADDRREADYTOACCEPT : in std_ulogic;
      MCMIREADDATA         : in std_logic_vector(0 to 127);
      MCMIREADDATAERR      : in std_ulogic;
      MCMIREADDATAVALID    : in std_ulogic;
      PLBPPCMADDRACK       : in std_ulogic;
      PLBPPCMMBUSY         : in std_ulogic;
      PLBPPCMMIRQ          : in std_ulogic;
      PLBPPCMMRDERR        : in std_ulogic;
      PLBPPCMMWRERR        : in std_ulogic;
      PLBPPCMRDBTERM       : in std_ulogic;
      PLBPPCMRDDACK        : in std_ulogic;
      PLBPPCMRDDBUS        : in std_logic_vector(0 to 127);
      PLBPPCMRDPENDPRI     : in std_logic_vector(0 to 1);
      PLBPPCMRDPENDREQ     : in std_ulogic;
      PLBPPCMRDWDADDR      : in std_logic_vector(0 to 3);
      PLBPPCMREARBITRATE   : in std_ulogic;
      PLBPPCMREQPRI        : in std_logic_vector(0 to 1);
      PLBPPCMSSIZE         : in std_logic_vector(0 to 1);
      PLBPPCMTIMEOUT       : in std_ulogic;
      PLBPPCMWRBTERM       : in std_ulogic;
      PLBPPCMWRDACK        : in std_ulogic;
      PLBPPCMWRPENDPRI     : in std_logic_vector(0 to 1);
      PLBPPCMWRPENDREQ     : in std_ulogic;
      PLBPPCS0ABORT        : in std_ulogic;
      PLBPPCS0ABUS         : in std_logic_vector(0 to 31);
      PLBPPCS0BE           : in std_logic_vector(0 to 15);
      PLBPPCS0BUSLOCK      : in std_ulogic;
      PLBPPCS0LOCKERR      : in std_ulogic;
      PLBPPCS0MASTERID     : in std_logic_vector(0 to 1);
      PLBPPCS0MSIZE        : in std_logic_vector(0 to 1);
      PLBPPCS0PAVALID      : in std_ulogic;
      PLBPPCS0RDBURST      : in std_ulogic;
      PLBPPCS0RDPENDPRI    : in std_logic_vector(0 to 1);
      PLBPPCS0RDPENDREQ    : in std_ulogic;
      PLBPPCS0RDPRIM       : in std_ulogic;
      PLBPPCS0REQPRI       : in std_logic_vector(0 to 1);
      PLBPPCS0RNW          : in std_ulogic;
      PLBPPCS0SAVALID      : in std_ulogic;
      PLBPPCS0SIZE         : in std_logic_vector(0 to 3);
      PLBPPCS0TATTRIBUTE   : in std_logic_vector(0 to 15);
      PLBPPCS0TYPE         : in std_logic_vector(0 to 2);
      PLBPPCS0UABUS        : in std_logic_vector(28 to 31);
      PLBPPCS0WRBURST      : in std_ulogic;
      PLBPPCS0WRDBUS       : in std_logic_vector(0 to 127);
      PLBPPCS0WRPENDPRI    : in std_logic_vector(0 to 1);
      PLBPPCS0WRPENDREQ    : in std_ulogic;
      PLBPPCS0WRPRIM       : in std_ulogic;
      PLBPPCS1ABORT        : in std_ulogic;
      PLBPPCS1ABUS         : in std_logic_vector(0 to 31);
      PLBPPCS1BE           : in std_logic_vector(0 to 15);
      PLBPPCS1BUSLOCK      : in std_ulogic;
      PLBPPCS1LOCKERR      : in std_ulogic;
      PLBPPCS1MASTERID     : in std_logic_vector(0 to 1);
      PLBPPCS1MSIZE        : in std_logic_vector(0 to 1);
      PLBPPCS1PAVALID      : in std_ulogic;
      PLBPPCS1RDBURST      : in std_ulogic;
      PLBPPCS1RDPENDPRI    : in std_logic_vector(0 to 1);
      PLBPPCS1RDPENDREQ    : in std_ulogic;
      PLBPPCS1RDPRIM       : in std_ulogic;
      PLBPPCS1REQPRI       : in std_logic_vector(0 to 1);
      PLBPPCS1RNW          : in std_ulogic;
      PLBPPCS1SAVALID      : in std_ulogic;
      PLBPPCS1SIZE         : in std_logic_vector(0 to 3);
      PLBPPCS1TATTRIBUTE   : in std_logic_vector(0 to 15);
      PLBPPCS1TYPE         : in std_logic_vector(0 to 2);
      PLBPPCS1UABUS        : in std_logic_vector(28 to 31);
      PLBPPCS1WRBURST      : in std_ulogic;
      PLBPPCS1WRDBUS       : in std_logic_vector(0 to 127);
      PLBPPCS1WRPENDPRI    : in std_logic_vector(0 to 1);
      PLBPPCS1WRPENDREQ    : in std_ulogic;
      PLBPPCS1WRPRIM       : in std_ulogic;
      RSTC440RESETCHIP     : in std_ulogic;
      RSTC440RESETCORE     : in std_ulogic;
      RSTC440RESETSYSTEM   : in std_ulogic;
      TIEC440DCURDLDCACHEPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440DCURDNONCACHEPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440DCURDTOUCHPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440DCURDURGENTPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440DCUWRFLUSHPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440DCUWRSTOREPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440DCUWRURGENTPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440ENDIANRESET   : in std_ulogic;
      TIEC440ERPNRESET     : in std_logic_vector(0 to 3);
      TIEC440ICURDFETCHPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440ICURDSPECPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440ICURDTOUCHPLBPRIO : in std_logic_vector(0 to 1);
      TIEC440PIR           : in std_logic_vector(28 to 31);
      TIEC440PVR           : in std_logic_vector(28 to 31);
      TIEC440USERRESET     : in std_logic_vector(0 to 3);
      TIEDCRBASEADDR       : in std_logic_vector(0 to 1);
      TRCC440TRACEDISABLE  : in std_ulogic;
      TRCC440TRIGGEREVENTIN : in std_ulogic;

      APU_CONTROL               : in std_logic_vector(0 to 16);
      APU_UDI0                  : in std_logic_vector(0 to 23);
      APU_UDI1                  : in std_logic_vector(0 to 23);
      APU_UDI10                 : in std_logic_vector(0 to 23);
      APU_UDI11                 : in std_logic_vector(0 to 23);
      APU_UDI12                 : in std_logic_vector(0 to 23);
      APU_UDI13                 : in std_logic_vector(0 to 23);
      APU_UDI14                 : in std_logic_vector(0 to 23);
      APU_UDI15                 : in std_logic_vector(0 to 23);
      APU_UDI2                  : in std_logic_vector(0 to 23);
      APU_UDI3                  : in std_logic_vector(0 to 23);
      APU_UDI4                  : in std_logic_vector(0 to 23);
      APU_UDI5                  : in std_logic_vector(0 to 23);
      APU_UDI6                  : in std_logic_vector(0 to 23);
      APU_UDI7                  : in std_logic_vector(0 to 23);
      APU_UDI8                  : in std_logic_vector(0 to 23);
      APU_UDI9                  : in std_logic_vector(0 to 23);
--      CLOCK_DELAY               : in std_ulogic;
      CLOCK_DELAY               : in std_logic_vector(0 to 4);
      DCR_AUTOLOCK_ENABLE       : in std_ulogic;
      DMA0_CONTROL              : in std_logic_vector(0 to 7);
      DMA0_RXCHANNELCTRL        : in std_logic_vector(0 to 31);
      DMA0_RXIRQTIMER           : in std_logic_vector(0 to 9);
      DMA0_TXCHANNELCTRL        : in std_logic_vector(0 to 31);
      DMA0_TXIRQTIMER           : in std_logic_vector(0 to 9);
      DMA1_CONTROL              : in std_logic_vector(0 to 7);
      DMA1_RXCHANNELCTRL        : in std_logic_vector(0 to 31);
      DMA1_RXIRQTIMER           : in std_logic_vector(0 to 9);
      DMA1_TXCHANNELCTRL        : in std_logic_vector(0 to 31);
      DMA1_TXIRQTIMER           : in std_logic_vector(0 to 9);
      DMA2_CONTROL              : in std_logic_vector(0 to 7);
      DMA2_RXCHANNELCTRL        : in std_logic_vector(0 to 31);
      DMA2_RXIRQTIMER           : in std_logic_vector(0 to 9);
      DMA2_TXCHANNELCTRL        : in std_logic_vector(0 to 31);
      DMA2_TXIRQTIMER           : in std_logic_vector(0 to 9);
      DMA3_CONTROL              : in std_logic_vector(0 to 7);
      DMA3_RXCHANNELCTRL        : in std_logic_vector(0 to 31);
      DMA3_RXIRQTIMER           : in std_logic_vector(0 to 9);
      DMA3_TXCHANNELCTRL        : in std_logic_vector(0 to 31);
      DMA3_TXIRQTIMER           : in std_logic_vector(0 to 9);
      INTERCONNECT_IMASK        : in std_logic_vector(0 to 31);
      INTERCONNECT_TMPL_SEL     : in std_logic_vector(0 to 31);
      MI_ARBCONFIG              : in std_logic_vector(0 to 31);
      MI_BANKCONFLICT_MASK      : in std_logic_vector(0 to 31);
      MI_CONTROL                : in std_logic_vector(0 to 31);
      MI_ROWCONFLICT_MASK       : in std_logic_vector(0 to 31);

      PPCDM_ASYNCMODE           : in std_ulogic;
      PPCDS_ASYNCMODE           : in std_ulogic;
      PPCM_ARBCONFIG            : in std_logic_vector(0 to 31);
      PPCM_CONTROL              : in std_logic_vector(0 to 31);
      PPCM_COUNTER              : in std_logic_vector(0 to 31);
      PPCS0_ADDRMAP_TMPL0       : in std_logic_vector(0 to 31);
      PPCS0_ADDRMAP_TMPL1       : in std_logic_vector(0 to 31);
      PPCS0_ADDRMAP_TMPL2       : in std_logic_vector(0 to 31);
      PPCS0_ADDRMAP_TMPL3       : in std_logic_vector(0 to 31);
      PPCS0_CONTROL             : in std_logic_vector(0 to 31);
      PPCS0_WIDTH_128N64        : in std_ulogic;
      PPCS1_ADDRMAP_TMPL0       : in std_logic_vector(0 to 31);
      PPCS1_ADDRMAP_TMPL1       : in std_logic_vector(0 to 31);
      PPCS1_ADDRMAP_TMPL2       : in std_logic_vector(0 to 31);
      PPCS1_ADDRMAP_TMPL3       : in std_logic_vector(0 to 31);
      PPCS1_CONTROL             : in std_logic_vector(0 to 31);
      PPCS1_WIDTH_128N64        : in std_ulogic;
      XBAR_ADDRMAP_TMPL0        : in std_logic_vector(0 to 31);
      XBAR_ADDRMAP_TMPL1        : in std_logic_vector(0 to 31);
      XBAR_ADDRMAP_TMPL2        : in std_logic_vector(0 to 31);
      XBAR_ADDRMAP_TMPL3        : in std_logic_vector(0 to 31)
    );
  end component;

	constant IN_DELAY : time :=  1 ps;
	constant OUT_DELAY : time := 0 ps;
	constant CLK_DELAY : time := 0 ps;

	signal   DMA3_TXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA3_TXCHANNELCTRL);
	signal   DMA3_CONTROL_BINARY  :  std_logic_vector(0 to 7) := To_StdLogicVector(DMA3_CONTROL);
	signal   DMA3_RXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA3_RXCHANNELCTRL);
	signal   DMA3_TXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA3_TXIRQTIMER)(9 downto 0);
	signal   DMA3_RXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA3_RXIRQTIMER)(9 downto 0);
	signal   DMA2_TXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA2_TXCHANNELCTRL);
	signal   DMA2_CONTROL_BINARY  :  std_logic_vector(0 to 7) := To_StdLogicVector(DMA2_CONTROL);
	signal   DMA2_RXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA2_RXCHANNELCTRL);
	signal   DMA2_TXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA2_TXIRQTIMER)(9 downto 0);
	signal   DMA2_RXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA2_RXIRQTIMER)(9 downto 0);
	signal   PPCM_CONTROL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCM_CONTROL);
	signal   PPCM_COUNTER_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCM_COUNTER);
	signal   PPCM_ARBCONFIG_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCM_ARBCONFIG);
	signal   DMA1_RXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA1_RXIRQTIMER)(9 downto 0);
	signal   DMA1_TXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA1_TXIRQTIMER)(9 downto 0);
	signal   DMA1_RXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA1_RXCHANNELCTRL);
	signal   DMA1_CONTROL_BINARY  :  std_logic_vector(0 to 7) := To_StdLogicVector(DMA1_CONTROL);
	signal   DMA1_TXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA1_TXCHANNELCTRL);
	signal   DMA0_RXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA0_RXIRQTIMER)(9 downto 0);
	signal   DMA0_TXIRQTIMER_BINARY  :  std_logic_vector(0 to 9) := To_StdLogicVector(DMA0_TXIRQTIMER)(9 downto 0);
	signal   DMA0_RXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA0_RXCHANNELCTRL);
	signal   DMA0_CONTROL_BINARY  :  std_logic_vector(0 to 7) := To_StdLogicVector(DMA0_CONTROL);
	signal   DMA0_TXCHANNELCTRL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(DMA0_TXCHANNELCTRL);
	signal   MI_ROWCONFLICT_MASK_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(MI_ROWCONFLICT_MASK);
	signal   MI_BANKCONFLICT_MASK_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(MI_BANKCONFLICT_MASK);
	signal   MI_ARBCONFIG_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(MI_ARBCONFIG);
	signal   MI_CONTROL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(MI_CONTROL);
	signal   APU_UDI0_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI0);
	signal   APU_UDI1_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI1);
	signal   APU_UDI2_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI2);
	signal   APU_UDI3_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI3);
	signal   APU_UDI4_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI4);
	signal   APU_UDI5_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI5);
	signal   APU_UDI6_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI6);
	signal   APU_UDI7_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI7);
	signal   APU_UDI8_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI8);
	signal   APU_UDI9_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI9);
	signal   APU_UDI10_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI10);
	signal   APU_UDI11_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI11);
	signal   APU_UDI12_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI12);
	signal   APU_UDI13_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI13);
	signal   APU_UDI14_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI14);
	signal   APU_UDI15_BINARY  :  std_logic_vector(0 to 23) := To_StdLogicVector(APU_UDI15);
	signal   APU_CONTROL_BINARY  :  std_logic_vector(0 to 16) := To_StdLogicVector(APU_CONTROL)(16 downto 0);
	signal   INTERCONNECT_IMASK_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(INTERCONNECT_IMASK);
	signal   XBAR_ADDRMAP_TMPL0_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(XBAR_ADDRMAP_TMPL0);
	signal   XBAR_ADDRMAP_TMPL1_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(XBAR_ADDRMAP_TMPL1);
	signal   XBAR_ADDRMAP_TMPL2_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(XBAR_ADDRMAP_TMPL2);
	signal   XBAR_ADDRMAP_TMPL3_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(XBAR_ADDRMAP_TMPL3);
	signal   INTERCONNECT_TMPL_SEL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(INTERCONNECT_TMPL_SEL);
	signal   PPCS0_CONTROL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS0_CONTROL);
	signal   PPCS0_WIDTH_128N64_BINARY  :  std_ulogic;
	signal   PPCS0_ADDRMAP_TMPL0_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS0_ADDRMAP_TMPL0);
	signal   PPCS0_ADDRMAP_TMPL1_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS0_ADDRMAP_TMPL1);
	signal   PPCS0_ADDRMAP_TMPL2_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS0_ADDRMAP_TMPL2);
	signal   PPCS0_ADDRMAP_TMPL3_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS0_ADDRMAP_TMPL3);
	signal   PPCS1_CONTROL_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS1_CONTROL);
	signal   PPCS1_WIDTH_128N64_BINARY  :  std_ulogic;
	signal   PPCS1_ADDRMAP_TMPL0_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS1_ADDRMAP_TMPL0);
	signal   PPCS1_ADDRMAP_TMPL1_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS1_ADDRMAP_TMPL1);
	signal   PPCS1_ADDRMAP_TMPL2_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS1_ADDRMAP_TMPL2);
	signal   PPCS1_ADDRMAP_TMPL3_BINARY  :  std_logic_vector(0 to 31) := To_StdLogicVector(PPCS1_ADDRMAP_TMPL3);
	signal   PPCDM_ASYNCMODE_BINARY  :  std_ulogic;
	signal   PPCDS_ASYNCMODE_BINARY  :  std_ulogic;
	signal   DCR_AUTOLOCK_ENABLE_BINARY  :  std_ulogic;
	signal   CLOCK_DELAY_BINARY  :   std_logic_vector(0 to 4);

	signal   DMA0LLRSTENGINEACK_out  :  std_ulogic;
	signal   DMA0LLRXDSTRDYN_out  :  std_ulogic;
	signal   DMA0LLTXD_out  :  std_logic_vector(0 to 31);
	signal   DMA0LLTXEOFN_out  :  std_ulogic;
	signal   DMA0LLTXEOPN_out  :  std_ulogic;
	signal   DMA0LLTXREM_out  :  std_logic_vector(0 to 3);
	signal   DMA0LLTXSOFN_out  :  std_ulogic;
	signal   DMA0LLTXSOPN_out  :  std_ulogic;
	signal   DMA0LLTXSRCRDYN_out  :  std_ulogic;
	signal   DMA0RXIRQ_out  :  std_ulogic;
	signal   DMA0TXIRQ_out  :  std_ulogic;
	signal   DMA1LLRSTENGINEACK_out  :  std_ulogic;
	signal   DMA1LLRXDSTRDYN_out  :  std_ulogic;
	signal   DMA1LLTXD_out  :  std_logic_vector(0 to 31);
	signal   DMA1LLTXEOFN_out  :  std_ulogic;
	signal   DMA1LLTXEOPN_out  :  std_ulogic;
	signal   DMA1LLTXREM_out  :  std_logic_vector(0 to 3);
	signal   DMA1LLTXSOFN_out  :  std_ulogic;
	signal   DMA1LLTXSOPN_out  :  std_ulogic;
	signal   DMA1LLTXSRCRDYN_out  :  std_ulogic;
	signal   DMA1RXIRQ_out  :  std_ulogic;
	signal   DMA1TXIRQ_out  :  std_ulogic;
	signal   DMA2LLRSTENGINEACK_out  :  std_ulogic;
	signal   DMA2LLRXDSTRDYN_out  :  std_ulogic;
	signal   DMA2LLTXD_out  :  std_logic_vector(0 to 31);
	signal   DMA2LLTXEOFN_out  :  std_ulogic;
	signal   DMA2LLTXEOPN_out  :  std_ulogic;
	signal   DMA2LLTXREM_out  :  std_logic_vector(0 to 3);
	signal   DMA2LLTXSOFN_out  :  std_ulogic;
	signal   DMA2LLTXSOPN_out  :  std_ulogic;
	signal   DMA2LLTXSRCRDYN_out  :  std_ulogic;
	signal   DMA2RXIRQ_out  :  std_ulogic;
	signal   DMA2TXIRQ_out  :  std_ulogic;
	signal   DMA3LLRSTENGINEACK_out  :  std_ulogic;
	signal   DMA3LLRXDSTRDYN_out  :  std_ulogic;
	signal   DMA3LLTXD_out  :  std_logic_vector(0 to 31);
	signal   DMA3LLTXEOFN_out  :  std_ulogic;
	signal   DMA3LLTXEOPN_out  :  std_ulogic;
	signal   DMA3LLTXREM_out  :  std_logic_vector(0 to 3);
	signal   DMA3LLTXSOFN_out  :  std_ulogic;
	signal   DMA3LLTXSOPN_out  :  std_ulogic;
	signal   DMA3LLTXSRCRDYN_out  :  std_ulogic;
	signal   DMA3RXIRQ_out  :  std_ulogic;
	signal   DMA3TXIRQ_out  :  std_ulogic;
	signal   PPCDMDCRABUS_out  :  std_logic_vector(0 to 9);
	signal   PPCDMDCRDBUSOUT_out  :  std_logic_vector(0 to 31);
	signal   PPCDMDCRREAD_out  :  std_ulogic;
	signal   PPCDMDCRUABUS_out  :  std_logic_vector(20 to 21);
	signal   PPCDMDCRWRITE_out  :  std_ulogic;
	signal   PPCMPLBABORT_out  :  std_ulogic;
	signal   PPCMPLBABUS_out  :  std_logic_vector(0 to 31);
	signal   PPCMPLBBE_out  :  std_logic_vector(0 to 15);
	signal   PPCMPLBBUSLOCK_out  :  std_ulogic;
	signal   PPCMPLBLOCKERR_out  :  std_ulogic;
	signal   PPCMPLBPRIORITY_out  :  std_logic_vector(0 to 1);
	signal   PPCMPLBRDBURST_out  :  std_ulogic;
	signal   PPCMPLBREQUEST_out  :  std_ulogic;
	signal   PPCMPLBRNW_out  :  std_ulogic;
	signal   PPCMPLBSIZE_out  :  std_logic_vector(0 to 3);
	signal   PPCMPLBTATTRIBUTE_out  :  std_logic_vector(0 to 15);
	signal   PPCMPLBTYPE_out  :  std_logic_vector(0 to 2);
	signal   PPCMPLBUABUS_out  :  std_logic_vector(28 to 31);
	signal   PPCMPLBWRBURST_out  :  std_ulogic;
	signal   PPCMPLBWRDBUS_out  :  std_logic_vector(0 to 127);
	signal   PPCS0PLBADDRACK_out  :  std_ulogic;
	signal   PPCS0PLBMBUSY_out  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBMIRQ_out  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBMRDERR_out  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBMWRERR_out  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBRDBTERM_out  :  std_ulogic;
	signal   PPCS0PLBRDCOMP_out  :  std_ulogic;
	signal   PPCS0PLBRDDACK_out  :  std_ulogic;
	signal   PPCS0PLBRDDBUS_out  :  std_logic_vector(0 to 127);
	signal   PPCS0PLBRDWDADDR_out  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBREARBITRATE_out  :  std_ulogic;
	signal   PPCS0PLBSSIZE_out  :  std_logic_vector(0 to 1);
	signal   PPCS0PLBWAIT_out  :  std_ulogic;
	signal   PPCS0PLBWRBTERM_out  :  std_ulogic;
	signal   PPCS0PLBWRCOMP_out  :  std_ulogic;
	signal   PPCS0PLBWRDACK_out  :  std_ulogic;
	signal   PPCS1PLBADDRACK_out  :  std_ulogic;
	signal   PPCS1PLBMBUSY_out  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBMIRQ_out  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBMRDERR_out  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBMWRERR_out  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBRDBTERM_out  :  std_ulogic;
	signal   PPCS1PLBRDCOMP_out  :  std_ulogic;
	signal   PPCS1PLBRDDACK_out  :  std_ulogic;
	signal   PPCS1PLBRDDBUS_out  :  std_logic_vector(0 to 127);
	signal   PPCS1PLBRDWDADDR_out  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBREARBITRATE_out  :  std_ulogic;
	signal   PPCS1PLBSSIZE_out  :  std_logic_vector(0 to 1);
	signal   PPCS1PLBWAIT_out  :  std_ulogic;
	signal   PPCS1PLBWRBTERM_out  :  std_ulogic;
	signal   PPCS1PLBWRCOMP_out  :  std_ulogic;
	signal   PPCS1PLBWRDACK_out  :  std_ulogic;
	signal   APUFCMDECFPUOP_out  :  std_ulogic;
	signal   APUFCMDECLDSTXFERSIZE_out  :  std_logic_vector(0 to 2);
	signal   APUFCMDECLOAD_out  :  std_ulogic;
	signal   APUFCMDECNONAUTON_out  :  std_ulogic;
	signal   APUFCMDECSTORE_out  :  std_ulogic;
	signal   APUFCMDECUDI_out  :  std_logic_vector(0 to 3);
	signal   APUFCMDECUDIVALID_out  :  std_ulogic;
	signal   APUFCMENDIAN_out  :  std_ulogic;
	signal   APUFCMFLUSH_out  :  std_ulogic;
	signal   APUFCMINSTRUCTION_out  :  std_logic_vector(0 to 31);
	signal   APUFCMINSTRVALID_out  :  std_ulogic;
	signal   APUFCMLOADBYTEADDR_out  :  std_logic_vector(0 to 3);
	signal   APUFCMLOADDATA_out  :  std_logic_vector(0 to 127);
	signal   APUFCMLOADDVALID_out  :  std_ulogic;
	signal   APUFCMMSRFE0_out  :  std_ulogic;
	signal   APUFCMMSRFE1_out  :  std_ulogic;
	signal   APUFCMNEXTINSTRREADY_out  :  std_ulogic;
	signal   APUFCMOPERANDVALID_out  :  std_ulogic;
	signal   APUFCMRADATA_out  :  std_logic_vector(0 to 31);
	signal   APUFCMRBDATA_out  :  std_logic_vector(0 to 31);
	signal   APUFCMWRITEBACKOK_out  :  std_ulogic;
	signal   C440CPMCORESLEEPREQ_out  :  std_ulogic;
	signal   C440CPMDECIRPTREQ_out  :  std_ulogic;
	signal   C440CPMFITIRPTREQ_out  :  std_ulogic;
	signal   C440CPMMSRCE_out  :  std_ulogic;
	signal   C440CPMMSREE_out  :  std_ulogic;
	signal   C440CPMTIMERRESETREQ_out  :  std_ulogic;
	signal   C440CPMWDIRPTREQ_out  :  std_ulogic;
	signal   C440DBGSYSTEMCONTROL_out  :  std_logic_vector(0 to 7);
	signal   C440JTGTDO_out  :  std_ulogic;
	signal   C440JTGTDOEN_out  :  std_ulogic;
	signal   C440MACHINECHECK_out  :  std_ulogic;
	signal   C440RSTCHIPRESETREQ_out  :  std_ulogic;
	signal   C440RSTCORERESETREQ_out  :  std_ulogic;
	signal   C440RSTSYSTEMRESETREQ_out  :  std_ulogic;
	signal   C440TRCBRANCHSTATUS_out  :  std_logic_vector(0 to 2);
	signal   C440TRCCYCLE_out  :  std_ulogic;
	signal   C440TRCEXECUTIONSTATUS_out  :  std_logic_vector(0 to 4);
	signal   C440TRCTRACESTATUS_out  :  std_logic_vector(0 to 6);
	signal   C440TRCTRIGGEREVENTOUT_out  :  std_ulogic;
	signal   C440TRCTRIGGEREVENTTYPE_out  :  std_logic_vector(0 to 13);
	signal   MIMCADDRESS_out  :  std_logic_vector(0 to 35);
	signal   MIMCADDRESSVALID_out  :  std_ulogic;
	signal   MIMCBANKCONFLICT_out  :  std_ulogic;
	signal   MIMCBYTEENABLE_out  :  std_logic_vector(0 to 15);
	signal   MIMCREADNOTWRITE_out  :  std_ulogic;
	signal   MIMCROWCONFLICT_out  :  std_ulogic;
	signal   MIMCWRITEDATA_out  :  std_logic_vector(0 to 127);
	signal   MIMCWRITEDATAVALID_out  :  std_ulogic;
	signal   PPCCPMINTERCONNECTBUSY_out  :  std_ulogic;
	signal   PPCDSDCRACK_out  :  std_ulogic;
	signal   PPCDSDCRTIMEOUTWAIT_out  :  std_ulogic;
	signal   PPCDSDCRDBUSIN_out  :  std_logic_vector(0 to 31);
	signal   PPCEICINTERCONNECTIRQ_out  :  std_ulogic;

	signal   DMA0LLRSTENGINEACK_outdelay  :  std_ulogic;
	signal   DMA0LLRXDSTRDYN_outdelay  :  std_ulogic;
	signal   DMA0LLTXD_outdelay  :  std_logic_vector(0 to 31);
	signal   DMA0LLTXEOFN_outdelay  :  std_ulogic;
	signal   DMA0LLTXEOPN_outdelay  :  std_ulogic;
	signal   DMA0LLTXREM_outdelay  :  std_logic_vector(0 to 3);
	signal   DMA0LLTXSOFN_outdelay  :  std_ulogic;
	signal   DMA0LLTXSOPN_outdelay  :  std_ulogic;
	signal   DMA0LLTXSRCRDYN_outdelay  :  std_ulogic;
	signal   DMA0RXIRQ_outdelay  :  std_ulogic;
	signal   DMA0TXIRQ_outdelay  :  std_ulogic;
	signal   DMA1LLRSTENGINEACK_outdelay  :  std_ulogic;
	signal   DMA1LLRXDSTRDYN_outdelay  :  std_ulogic;
	signal   DMA1LLTXD_outdelay  :  std_logic_vector(0 to 31);
	signal   DMA1LLTXEOFN_outdelay  :  std_ulogic;
	signal   DMA1LLTXEOPN_outdelay  :  std_ulogic;
	signal   DMA1LLTXREM_outdelay  :  std_logic_vector(0 to 3);
	signal   DMA1LLTXSOFN_outdelay  :  std_ulogic;
	signal   DMA1LLTXSOPN_outdelay  :  std_ulogic;
	signal   DMA1LLTXSRCRDYN_outdelay  :  std_ulogic;
	signal   DMA1RXIRQ_outdelay  :  std_ulogic;
	signal   DMA1TXIRQ_outdelay  :  std_ulogic;
	signal   DMA2LLRSTENGINEACK_outdelay  :  std_ulogic;
	signal   DMA2LLRXDSTRDYN_outdelay  :  std_ulogic;
	signal   DMA2LLTXD_outdelay  :  std_logic_vector(0 to 31);
	signal   DMA2LLTXEOFN_outdelay  :  std_ulogic;
	signal   DMA2LLTXEOPN_outdelay  :  std_ulogic;
	signal   DMA2LLTXREM_outdelay  :  std_logic_vector(0 to 3);
	signal   DMA2LLTXSOFN_outdelay  :  std_ulogic;
	signal   DMA2LLTXSOPN_outdelay  :  std_ulogic;
	signal   DMA2LLTXSRCRDYN_outdelay  :  std_ulogic;
	signal   DMA2RXIRQ_outdelay  :  std_ulogic;
	signal   DMA2TXIRQ_outdelay  :  std_ulogic;
	signal   DMA3LLRSTENGINEACK_outdelay  :  std_ulogic;
	signal   DMA3LLRXDSTRDYN_outdelay  :  std_ulogic;
	signal   DMA3LLTXD_outdelay  :  std_logic_vector(0 to 31);
	signal   DMA3LLTXEOFN_outdelay  :  std_ulogic;
	signal   DMA3LLTXEOPN_outdelay  :  std_ulogic;
	signal   DMA3LLTXREM_outdelay  :  std_logic_vector(0 to 3);
	signal   DMA3LLTXSOFN_outdelay  :  std_ulogic;
	signal   DMA3LLTXSOPN_outdelay  :  std_ulogic;
	signal   DMA3LLTXSRCRDYN_outdelay  :  std_ulogic;
	signal   DMA3RXIRQ_outdelay  :  std_ulogic;
	signal   DMA3TXIRQ_outdelay  :  std_ulogic;
	signal   PPCDMDCRABUS_outdelay  :  std_logic_vector(0 to 9);
	signal   PPCDMDCRDBUSOUT_outdelay  :  std_logic_vector(0 to 31);
	signal   PPCDMDCRREAD_outdelay  :  std_ulogic;
	signal   PPCDMDCRUABUS_outdelay  :  std_logic_vector(20 to 21);
	signal   PPCDMDCRWRITE_outdelay  :  std_ulogic;
	signal   PPCMPLBABORT_outdelay  :  std_ulogic;
	signal   PPCMPLBABUS_outdelay  :  std_logic_vector(0 to 31);
	signal   PPCMPLBBE_outdelay  :  std_logic_vector(0 to 15);
	signal   PPCMPLBBUSLOCK_outdelay  :  std_ulogic;
	signal   PPCMPLBLOCKERR_outdelay  :  std_ulogic;
	signal   PPCMPLBPRIORITY_outdelay  :  std_logic_vector(0 to 1);
	signal   PPCMPLBRDBURST_outdelay  :  std_ulogic;
	signal   PPCMPLBREQUEST_outdelay  :  std_ulogic;
	signal   PPCMPLBRNW_outdelay  :  std_ulogic;
	signal   PPCMPLBSIZE_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCMPLBTATTRIBUTE_outdelay  :  std_logic_vector(0 to 15);
	signal   PPCMPLBTYPE_outdelay  :  std_logic_vector(0 to 2);
	signal   PPCMPLBUABUS_outdelay  :  std_logic_vector(28 to 31);
	signal   PPCMPLBWRBURST_outdelay  :  std_ulogic;
	signal   PPCMPLBWRDBUS_outdelay  :  std_logic_vector(0 to 127);
	signal   PPCS0PLBADDRACK_outdelay  :  std_ulogic;
	signal   PPCS0PLBMBUSY_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBMIRQ_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBMRDERR_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBMWRERR_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBRDBTERM_outdelay  :  std_ulogic;
	signal   PPCS0PLBRDCOMP_outdelay  :  std_ulogic;
	signal   PPCS0PLBRDDACK_outdelay  :  std_ulogic;
	signal   PPCS0PLBRDDBUS_outdelay  :  std_logic_vector(0 to 127);
	signal   PPCS0PLBRDWDADDR_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS0PLBREARBITRATE_outdelay  :  std_ulogic;
	signal   PPCS0PLBSSIZE_outdelay  :  std_logic_vector(0 to 1);
	signal   PPCS0PLBWAIT_outdelay  :  std_ulogic;
	signal   PPCS0PLBWRBTERM_outdelay  :  std_ulogic;
	signal   PPCS0PLBWRCOMP_outdelay  :  std_ulogic;
	signal   PPCS0PLBWRDACK_outdelay  :  std_ulogic;
	signal   PPCS1PLBADDRACK_outdelay  :  std_ulogic;
	signal   PPCS1PLBMBUSY_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBMIRQ_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBMRDERR_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBMWRERR_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBRDBTERM_outdelay  :  std_ulogic;
	signal   PPCS1PLBRDCOMP_outdelay  :  std_ulogic;
	signal   PPCS1PLBRDDACK_outdelay  :  std_ulogic;
	signal   PPCS1PLBRDDBUS_outdelay  :  std_logic_vector(0 to 127);
	signal   PPCS1PLBRDWDADDR_outdelay  :  std_logic_vector(0 to 3);
	signal   PPCS1PLBREARBITRATE_outdelay  :  std_ulogic;
	signal   PPCS1PLBSSIZE_outdelay  :  std_logic_vector(0 to 1);
	signal   PPCS1PLBWAIT_outdelay  :  std_ulogic;
	signal   PPCS1PLBWRBTERM_outdelay  :  std_ulogic;
	signal   PPCS1PLBWRCOMP_outdelay  :  std_ulogic;
	signal   PPCS1PLBWRDACK_outdelay  :  std_ulogic;
	signal   APUFCMDECFPUOP_outdelay  :  std_ulogic;
	signal   APUFCMDECLDSTXFERSIZE_outdelay  :  std_logic_vector(0 to 2);
	signal   APUFCMDECLOAD_outdelay  :  std_ulogic;
	signal   APUFCMDECNONAUTON_outdelay  :  std_ulogic;
	signal   APUFCMDECSTORE_outdelay  :  std_ulogic;
	signal   APUFCMDECUDI_outdelay  :  std_logic_vector(0 to 3);
	signal   APUFCMDECUDIVALID_outdelay  :  std_ulogic;
	signal   APUFCMENDIAN_outdelay  :  std_ulogic;
	signal   APUFCMFLUSH_outdelay  :  std_ulogic;
	signal   APUFCMINSTRUCTION_outdelay  :  std_logic_vector(0 to 31);
	signal   APUFCMINSTRVALID_outdelay  :  std_ulogic;
	signal   APUFCMLOADBYTEADDR_outdelay  :  std_logic_vector(0 to 3);
	signal   APUFCMLOADDATA_outdelay  :  std_logic_vector(0 to 127);
	signal   APUFCMLOADDVALID_outdelay  :  std_ulogic;
	signal   APUFCMMSRFE0_outdelay  :  std_ulogic;
	signal   APUFCMMSRFE1_outdelay  :  std_ulogic;
	signal   APUFCMNEXTINSTRREADY_outdelay  :  std_ulogic;
	signal   APUFCMOPERANDVALID_outdelay  :  std_ulogic;
	signal   APUFCMRADATA_outdelay  :  std_logic_vector(0 to 31);
	signal   APUFCMRBDATA_outdelay  :  std_logic_vector(0 to 31);
	signal   APUFCMWRITEBACKOK_outdelay  :  std_ulogic;
	signal   C440CPMCORESLEEPREQ_outdelay  :  std_ulogic;
	signal   C440CPMDECIRPTREQ_outdelay  :  std_ulogic;
	signal   C440CPMFITIRPTREQ_outdelay  :  std_ulogic;
	signal   C440CPMMSRCE_outdelay  :  std_ulogic;
	signal   C440CPMMSREE_outdelay  :  std_ulogic;
	signal   C440CPMTIMERRESETREQ_outdelay  :  std_ulogic;
	signal   C440CPMWDIRPTREQ_outdelay  :  std_ulogic;
	signal   C440DBGSYSTEMCONTROL_outdelay  :  std_logic_vector(0 to 7);
	signal   C440JTGTDO_outdelay  :  std_ulogic;
	signal   C440JTGTDOEN_outdelay  :  std_ulogic;
	signal   C440MACHINECHECK_outdelay  :  std_ulogic;
	signal   C440RSTCHIPRESETREQ_outdelay  :  std_ulogic;
	signal   C440RSTCORERESETREQ_outdelay  :  std_ulogic;
	signal   C440RSTSYSTEMRESETREQ_outdelay  :  std_ulogic;
	signal   C440TRCBRANCHSTATUS_outdelay  :  std_logic_vector(0 to 2);
	signal   C440TRCCYCLE_outdelay  :  std_ulogic;
	signal   C440TRCEXECUTIONSTATUS_outdelay  :  std_logic_vector(0 to 4);
	signal   C440TRCTRACESTATUS_outdelay  :  std_logic_vector(0 to 6);
	signal   C440TRCTRIGGEREVENTOUT_outdelay  :  std_ulogic;
	signal   C440TRCTRIGGEREVENTTYPE_outdelay  :  std_logic_vector(0 to 13);
	signal   MIMCADDRESS_outdelay  :  std_logic_vector(0 to 35);
	signal   MIMCADDRESSVALID_outdelay  :  std_ulogic;
	signal   MIMCBANKCONFLICT_outdelay  :  std_ulogic;
	signal   MIMCBYTEENABLE_outdelay  :  std_logic_vector(0 to 15);
	signal   MIMCREADNOTWRITE_outdelay  :  std_ulogic;
	signal   MIMCROWCONFLICT_outdelay  :  std_ulogic;
	signal   MIMCWRITEDATA_outdelay  :  std_logic_vector(0 to 127);
	signal   MIMCWRITEDATAVALID_outdelay  :  std_ulogic;
	signal   PPCCPMINTERCONNECTBUSY_outdelay  :  std_ulogic;
	signal   PPCDSDCRACK_outdelay  :  std_ulogic;
	signal   PPCDSDCRTIMEOUTWAIT_outdelay  :  std_ulogic;
	signal   PPCDSDCRDBUSIN_outdelay  :  std_logic_vector(0 to 31);
	signal   PPCEICINTERCONNECTIRQ_outdelay  :  std_ulogic;

	signal   PLBPPCS0RNW_ipd  :  std_ulogic;
	signal   PLBPPCS1RNW_ipd  :  std_ulogic;
	signal   CPMDCRCLK_ipd  :  std_ulogic;
	signal   CPMDMA0LLCLK_ipd  :  std_ulogic;
	signal   CPMDMA1LLCLK_ipd  :  std_ulogic;
	signal   CPMDMA2LLCLK_ipd  :  std_ulogic;
	signal   CPMDMA3LLCLK_ipd  :  std_ulogic;
	signal   CPMINTERCONNECTCLKNTO1_ipd  :  std_ulogic;
	signal   CPMPPCMPLBCLK_ipd  :  std_ulogic;
	signal   CPMPPCS0PLBCLK_ipd  :  std_ulogic;
	signal   CPMPPCS1PLBCLK_ipd  :  std_ulogic;
	signal   DCRPPCDMACK_ipd  :  std_ulogic;
	signal   DCRPPCDMDBUSIN_ipd  :  std_logic_vector(0 to 31);
	signal   DCRPPCDMTIMEOUTWAIT_ipd  :  std_ulogic;
	signal   LLDMA0RSTENGINEREQ_ipd  :  std_ulogic;
	signal   LLDMA0RXD_ipd  :  std_logic_vector(0 to 31);
	signal   LLDMA0RXEOFN_ipd  :  std_ulogic;
	signal   LLDMA0RXEOPN_ipd  :  std_ulogic;
	signal   LLDMA0RXREM_ipd  :  std_logic_vector(0 to 3);
	signal   LLDMA0RXSOFN_ipd  :  std_ulogic;
	signal   LLDMA0RXSOPN_ipd  :  std_ulogic;
	signal   LLDMA0RXSRCRDYN_ipd  :  std_ulogic;
	signal   LLDMA0TXDSTRDYN_ipd  :  std_ulogic;
	signal   LLDMA1RSTENGINEREQ_ipd  :  std_ulogic;
	signal   LLDMA1RXD_ipd  :  std_logic_vector(0 to 31);
	signal   LLDMA1RXEOFN_ipd  :  std_ulogic;
	signal   LLDMA1RXEOPN_ipd  :  std_ulogic;
	signal   LLDMA1RXREM_ipd  :  std_logic_vector(0 to 3);
	signal   LLDMA1RXSOFN_ipd  :  std_ulogic;
	signal   LLDMA1RXSOPN_ipd  :  std_ulogic;
	signal   LLDMA1RXSRCRDYN_ipd  :  std_ulogic;
	signal   LLDMA1TXDSTRDYN_ipd  :  std_ulogic;
	signal   LLDMA2RSTENGINEREQ_ipd  :  std_ulogic;
	signal   LLDMA2RXD_ipd  :  std_logic_vector(0 to 31);
	signal   LLDMA2RXEOFN_ipd  :  std_ulogic;
	signal   LLDMA2RXEOPN_ipd  :  std_ulogic;
	signal   LLDMA2RXREM_ipd  :  std_logic_vector(0 to 3);
	signal   LLDMA2RXSOFN_ipd  :  std_ulogic;
	signal   LLDMA2RXSOPN_ipd  :  std_ulogic;
	signal   LLDMA2RXSRCRDYN_ipd  :  std_ulogic;
	signal   LLDMA2TXDSTRDYN_ipd  :  std_ulogic;
	signal   LLDMA3RSTENGINEREQ_ipd  :  std_ulogic;
	signal   LLDMA3RXD_ipd  :  std_logic_vector(0 to 31);
	signal   LLDMA3RXEOFN_ipd  :  std_ulogic;
	signal   LLDMA3RXEOPN_ipd  :  std_ulogic;
	signal   LLDMA3RXREM_ipd  :  std_logic_vector(0 to 3);
	signal   LLDMA3RXSOFN_ipd  :  std_ulogic;
	signal   LLDMA3RXSOPN_ipd  :  std_ulogic;
	signal   LLDMA3RXSRCRDYN_ipd  :  std_ulogic;
	signal   LLDMA3TXDSTRDYN_ipd  :  std_ulogic;
	signal   PLBPPCMADDRACK_ipd  :  std_ulogic;
	signal   PLBPPCMMBUSY_ipd  :  std_ulogic;
	signal   PLBPPCMMIRQ_ipd  :  std_ulogic;
	signal   PLBPPCMMRDERR_ipd  :  std_ulogic;
	signal   PLBPPCMMWRERR_ipd  :  std_ulogic;
	signal   PLBPPCMRDBTERM_ipd  :  std_ulogic;
	signal   PLBPPCMRDDACK_ipd  :  std_ulogic;
	signal   PLBPPCMRDDBUS_ipd  :  std_logic_vector(0 to 127);
	signal   PLBPPCMRDPENDPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCMRDPENDREQ_ipd  :  std_ulogic;
	signal   PLBPPCMRDWDADDR_ipd  :  std_logic_vector(0 to 3);
	signal   PLBPPCMREARBITRATE_ipd  :  std_ulogic;
	signal   PLBPPCMREQPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCMSSIZE_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCMTIMEOUT_ipd  :  std_ulogic;
	signal   PLBPPCMWRBTERM_ipd  :  std_ulogic;
	signal   PLBPPCMWRDACK_ipd  :  std_ulogic;
	signal   PLBPPCMWRPENDPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCMWRPENDREQ_ipd  :  std_ulogic;
	signal   PLBPPCS0ABORT_ipd  :  std_ulogic;
	signal   PLBPPCS0ABUS_ipd  :  std_logic_vector(0 to 31);
	signal   PLBPPCS0BE_ipd  :  std_logic_vector(0 to 15);
	signal   PLBPPCS0BUSLOCK_ipd  :  std_ulogic;
	signal   PLBPPCS0LOCKERR_ipd  :  std_ulogic;
	signal   PLBPPCS0MASTERID_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0MSIZE_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0PAVALID_ipd  :  std_ulogic;
	signal   PLBPPCS0RDBURST_ipd  :  std_ulogic;
	signal   PLBPPCS0RDPENDPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0RDPENDREQ_ipd  :  std_ulogic;
	signal   PLBPPCS0RDPRIM_ipd  :  std_ulogic;
	signal   PLBPPCS0REQPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0SAVALID_ipd  :  std_ulogic;
	signal   PLBPPCS0SIZE_ipd  :  std_logic_vector(0 to 3);
	signal   PLBPPCS0TATTRIBUTE_ipd  :  std_logic_vector(0 to 15);
	signal   PLBPPCS0TYPE_ipd  :  std_logic_vector(0 to 2);
	signal   PLBPPCS0UABUS_ipd  :  std_logic_vector(28 to 31);
	signal   PLBPPCS0WRBURST_ipd  :  std_ulogic;
	signal   PLBPPCS0WRDBUS_ipd  :  std_logic_vector(0 to 127);
	signal   PLBPPCS0WRPENDPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0WRPENDREQ_ipd  :  std_ulogic;
	signal   PLBPPCS0WRPRIM_ipd  :  std_ulogic;
	signal   PLBPPCS1ABORT_ipd  :  std_ulogic;
	signal   PLBPPCS1ABUS_ipd  :  std_logic_vector(0 to 31);
	signal   PLBPPCS1BE_ipd  :  std_logic_vector(0 to 15);
	signal   PLBPPCS1BUSLOCK_ipd  :  std_ulogic;
	signal   PLBPPCS1LOCKERR_ipd  :  std_ulogic;
	signal   PLBPPCS1MASTERID_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1MSIZE_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1PAVALID_ipd  :  std_ulogic;
	signal   PLBPPCS1RDBURST_ipd  :  std_ulogic;
	signal   PLBPPCS1RDPENDPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1RDPENDREQ_ipd  :  std_ulogic;
	signal   PLBPPCS1RDPRIM_ipd  :  std_ulogic;
	signal   PLBPPCS1REQPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1SAVALID_ipd  :  std_ulogic;
	signal   PLBPPCS1SIZE_ipd  :  std_logic_vector(0 to 3);
	signal   PLBPPCS1TATTRIBUTE_ipd  :  std_logic_vector(0 to 15);
	signal   PLBPPCS1TYPE_ipd  :  std_logic_vector(0 to 2);
	signal   PLBPPCS1UABUS_ipd  :  std_logic_vector(28 to 31);
	signal   PLBPPCS1WRBURST_ipd  :  std_ulogic;
	signal   PLBPPCS1WRDBUS_ipd  :  std_logic_vector(0 to 127);
	signal   PLBPPCS1WRPENDPRI_ipd  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1WRPENDREQ_ipd  :  std_ulogic;
	signal   PLBPPCS1WRPRIM_ipd  :  std_ulogic;
	signal   TIEDCRBASEADDR_ipd  :  std_logic_vector(0 to 1);
	signal   CPMC440CLK_ipd  :  std_ulogic;
	signal   CPMC440CLKEN_ipd  :  std_ulogic;
	signal   CPMC440CORECLOCKINACTIVE_ipd  :  std_ulogic;
	signal   CPMC440TIMERCLOCK_ipd  :  std_ulogic;
	signal   CPMFCMCLK_ipd  :  std_ulogic;
	signal   CPMINTERCONNECTCLK_ipd  :  std_ulogic;
	signal   CPMINTERCONNECTCLKEN_ipd  :  std_ulogic;
	signal   CPMMCCLK_ipd  :  std_ulogic;
	signal   DBGC440DEBUGHALT_ipd  :  std_ulogic;
	signal   DBGC440SYSTEMSTATUS_ipd  :  std_logic_vector(0 to 4);
	signal   DBGC440UNCONDDEBUGEVENT_ipd  :  std_ulogic;
	signal   DCRPPCDSABUS_ipd  :  std_logic_vector(0 to 9);
	signal   DCRPPCDSDBUSOUT_ipd  :  std_logic_vector(0 to 31);
	signal   DCRPPCDSREAD_ipd  :  std_ulogic;
	signal   DCRPPCDSWRITE_ipd  :  std_ulogic;
	signal   EICC440CRITIRQ_ipd  :  std_ulogic;
	signal   EICC440EXTIRQ_ipd  :  std_ulogic;
	signal   FCMAPUCONFIRMINSTR_ipd  :  std_ulogic;
	signal   FCMAPUCR_ipd  :  std_logic_vector(0 to 3);
	signal   FCMAPUDONE_ipd  :  std_ulogic;
	signal   FCMAPUEXCEPTION_ipd  :  std_ulogic;
	signal   FCMAPUFPSCRFEX_ipd  :  std_ulogic;
	signal   FCMAPURESULT_ipd  :  std_logic_vector(0 to 31);
	signal   FCMAPURESULTVALID_ipd  :  std_ulogic;
	signal   FCMAPUSLEEPNOTREADY_ipd  :  std_ulogic;
	signal   FCMAPUSTOREDATA_ipd  :  std_logic_vector(0 to 127);
	signal   JTGC440TCK_ipd  :  std_ulogic;
	signal   JTGC440TDI_ipd  :  std_ulogic;
	signal   JTGC440TMS_ipd  :  std_ulogic;
	signal   JTGC440TRSTNEG_ipd  :  std_ulogic;
	signal   MCMIADDRREADYTOACCEPT_ipd  :  std_ulogic;
	signal   MCMIREADDATA_ipd  :  std_logic_vector(0 to 127);
	signal   MCMIREADDATAERR_ipd  :  std_ulogic;
	signal   MCMIREADDATAVALID_ipd  :  std_ulogic;
	signal   RSTC440RESETCHIP_ipd  :  std_ulogic;
	signal   RSTC440RESETCORE_ipd  :  std_ulogic;
	signal   RSTC440RESETSYSTEM_ipd  :  std_ulogic;
	signal   TIEC440DCURDLDCACHEPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDNONCACHEPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDTOUCHPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDURGENTPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRFLUSHPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRSTOREPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRURGENTPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440ENDIANRESET_ipd  :  std_ulogic;
	signal   TIEC440ERPNRESET_ipd  :  std_logic_vector(0 to 3);
	signal   TIEC440ICURDFETCHPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440ICURDSPECPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440ICURDTOUCHPLBPRIO_ipd  :  std_logic_vector(0 to 1);
	signal   TIEC440PIR_ipd  :  std_logic_vector(28 to 31);
	signal   TIEC440PVR_ipd  :  std_logic_vector(28 to 31);
	signal   TIEC440USERRESET_ipd  :  std_logic_vector(0 to 3);
	signal   TRCC440TRACEDISABLE_ipd  :  std_ulogic;
	signal   TRCC440TRIGGEREVENTIN_ipd  :  std_ulogic;

	signal   PLBPPCS0RNW_dly  :  std_ulogic;
	signal   PLBPPCS1RNW_dly  :  std_ulogic;
	signal   CPMDCRCLK_dly  :  std_ulogic;
	signal   CPMDMA0LLCLK_dly  :  std_ulogic;
	signal   CPMDMA1LLCLK_dly  :  std_ulogic;
	signal   CPMDMA2LLCLK_dly  :  std_ulogic;
	signal   CPMDMA3LLCLK_dly  :  std_ulogic;
	signal   CPMINTERCONNECTCLKNTO1_dly  :  std_ulogic;
	signal   CPMPPCMPLBCLK_dly  :  std_ulogic;
	signal   CPMPPCS0PLBCLK_dly  :  std_ulogic;
	signal   CPMPPCS1PLBCLK_dly  :  std_ulogic;
	signal   DCRPPCDMACK_dly  :  std_ulogic;
	signal   DCRPPCDMDBUSIN_dly  :  std_logic_vector(0 to 31);
	signal   DCRPPCDMTIMEOUTWAIT_dly  :  std_ulogic;
	signal   LLDMA0RSTENGINEREQ_dly  :  std_ulogic;
	signal   LLDMA0RXD_dly  :  std_logic_vector(0 to 31);
	signal   LLDMA0RXEOFN_dly  :  std_ulogic;
	signal   LLDMA0RXEOPN_dly  :  std_ulogic;
	signal   LLDMA0RXREM_dly  :  std_logic_vector(0 to 3);
	signal   LLDMA0RXSOFN_dly  :  std_ulogic;
	signal   LLDMA0RXSOPN_dly  :  std_ulogic;
	signal   LLDMA0RXSRCRDYN_dly  :  std_ulogic;
	signal   LLDMA0TXDSTRDYN_dly  :  std_ulogic;
	signal   LLDMA1RSTENGINEREQ_dly  :  std_ulogic;
	signal   LLDMA1RXD_dly  :  std_logic_vector(0 to 31);
	signal   LLDMA1RXEOFN_dly  :  std_ulogic;
	signal   LLDMA1RXEOPN_dly  :  std_ulogic;
	signal   LLDMA1RXREM_dly  :  std_logic_vector(0 to 3);
	signal   LLDMA1RXSOFN_dly  :  std_ulogic;
	signal   LLDMA1RXSOPN_dly  :  std_ulogic;
	signal   LLDMA1RXSRCRDYN_dly  :  std_ulogic;
	signal   LLDMA1TXDSTRDYN_dly  :  std_ulogic;
	signal   LLDMA2RSTENGINEREQ_dly  :  std_ulogic;
	signal   LLDMA2RXD_dly  :  std_logic_vector(0 to 31);
	signal   LLDMA2RXEOFN_dly  :  std_ulogic;
	signal   LLDMA2RXEOPN_dly  :  std_ulogic;
	signal   LLDMA2RXREM_dly  :  std_logic_vector(0 to 3);
	signal   LLDMA2RXSOFN_dly  :  std_ulogic;
	signal   LLDMA2RXSOPN_dly  :  std_ulogic;
	signal   LLDMA2RXSRCRDYN_dly  :  std_ulogic;
	signal   LLDMA2TXDSTRDYN_dly  :  std_ulogic;
	signal   LLDMA3RSTENGINEREQ_dly  :  std_ulogic;
	signal   LLDMA3RXD_dly  :  std_logic_vector(0 to 31);
	signal   LLDMA3RXEOFN_dly  :  std_ulogic;
	signal   LLDMA3RXEOPN_dly  :  std_ulogic;
	signal   LLDMA3RXREM_dly  :  std_logic_vector(0 to 3);
	signal   LLDMA3RXSOFN_dly  :  std_ulogic;
	signal   LLDMA3RXSOPN_dly  :  std_ulogic;
	signal   LLDMA3RXSRCRDYN_dly  :  std_ulogic;
	signal   LLDMA3TXDSTRDYN_dly  :  std_ulogic;
	signal   PLBPPCMADDRACK_dly  :  std_ulogic;
	signal   PLBPPCMMBUSY_dly  :  std_ulogic;
	signal   PLBPPCMMIRQ_dly  :  std_ulogic;
	signal   PLBPPCMMRDERR_dly  :  std_ulogic;
	signal   PLBPPCMMWRERR_dly  :  std_ulogic;
	signal   PLBPPCMRDBTERM_dly  :  std_ulogic;
	signal   PLBPPCMRDDACK_dly  :  std_ulogic;
	signal   PLBPPCMRDDBUS_dly  :  std_logic_vector(0 to 127);
	signal   PLBPPCMRDPENDPRI_dly  :  std_logic_vector(0 to 1);
	signal   PLBPPCMRDPENDREQ_dly  :  std_ulogic;
	signal   PLBPPCMRDWDADDR_dly  :  std_logic_vector(0 to 3);
	signal   PLBPPCMREARBITRATE_dly  :  std_ulogic;
	signal   PLBPPCMREQPRI_dly  :  std_logic_vector(0 to 1);
	signal   PLBPPCMSSIZE_dly  :  std_logic_vector(0 to 1);
	signal   PLBPPCMTIMEOUT_dly  :  std_ulogic;
	signal   PLBPPCMWRBTERM_dly  :  std_ulogic;
	signal   PLBPPCMWRDACK_dly  :  std_ulogic;
	signal   PLBPPCMWRPENDPRI_dly  :  std_logic_vector(0 to 1);
	signal   PLBPPCMWRPENDREQ_dly  :  std_ulogic;
	signal   PLBPPCS0ABORT_dly  :  std_ulogic;
	signal   PLBPPCS0ABUS_dly  :  std_logic_vector(0 to 31);
	signal   PLBPPCS0BE_dly  :  std_logic_vector(0 to 15);
	signal   PLBPPCS0BUSLOCK_dly  :  std_ulogic;
	signal   PLBPPCS0LOCKERR_dly  :  std_ulogic;
	signal   PLBPPCS0MASTERID_dly  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0MSIZE_dly  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0PAVALID_dly  :  std_ulogic;
	signal   PLBPPCS0RDBURST_dly  :  std_ulogic;
	signal   PLBPPCS0RDPENDPRI_dly  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0RDPENDREQ_dly  :  std_ulogic;
	signal   PLBPPCS0RDPRIM_dly  :  std_ulogic;
	signal   PLBPPCS0REQPRI_dly  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0SAVALID_dly  :  std_ulogic;
	signal   PLBPPCS0SIZE_dly  :  std_logic_vector(0 to 3);
	signal   PLBPPCS0TATTRIBUTE_dly  :  std_logic_vector(0 to 15);
	signal   PLBPPCS0TYPE_dly  :  std_logic_vector(0 to 2);
	signal   PLBPPCS0UABUS_dly  :  std_logic_vector(28 to 31);
	signal   PLBPPCS0WRBURST_dly  :  std_ulogic;
	signal   PLBPPCS0WRDBUS_dly  :  std_logic_vector(0 to 127);
	signal   PLBPPCS0WRPENDPRI_dly  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0WRPENDREQ_dly  :  std_ulogic;
	signal   PLBPPCS0WRPRIM_dly  :  std_ulogic;
	signal   PLBPPCS1ABORT_dly  :  std_ulogic;
	signal   PLBPPCS1ABUS_dly  :  std_logic_vector(0 to 31);
	signal   PLBPPCS1BE_dly  :  std_logic_vector(0 to 15);
	signal   PLBPPCS1BUSLOCK_dly  :  std_ulogic;
	signal   PLBPPCS1LOCKERR_dly  :  std_ulogic;
	signal   PLBPPCS1MASTERID_dly  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1MSIZE_dly  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1PAVALID_dly  :  std_ulogic;
	signal   PLBPPCS1RDBURST_dly  :  std_ulogic;
	signal   PLBPPCS1RDPENDPRI_dly  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1RDPENDREQ_dly  :  std_ulogic;
	signal   PLBPPCS1RDPRIM_dly  :  std_ulogic;
	signal   PLBPPCS1REQPRI_dly  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1SAVALID_dly  :  std_ulogic;
	signal   PLBPPCS1SIZE_dly  :  std_logic_vector(0 to 3);
	signal   PLBPPCS1TATTRIBUTE_dly  :  std_logic_vector(0 to 15);
	signal   PLBPPCS1TYPE_dly  :  std_logic_vector(0 to 2);
	signal   PLBPPCS1UABUS_dly  :  std_logic_vector(28 to 31);
	signal   PLBPPCS1WRBURST_dly  :  std_ulogic;
	signal   PLBPPCS1WRDBUS_dly  :  std_logic_vector(0 to 127);
	signal   PLBPPCS1WRPENDPRI_dly  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1WRPENDREQ_dly  :  std_ulogic;
	signal   PLBPPCS1WRPRIM_dly  :  std_ulogic;
	signal   TIEDCRBASEADDR_dly  :  std_logic_vector(0 to 1);
	signal   CPMC440CLK_dly  :  std_ulogic;
	signal   CPMC440CLKEN_dly  :  std_ulogic;
	signal   CPMC440CORECLOCKINACTIVE_dly  :  std_ulogic;
	signal   CPMC440TIMERCLOCK_dly  :  std_ulogic;
	signal   CPMFCMCLK_dly  :  std_ulogic;
	signal   CPMINTERCONNECTCLK_dly  :  std_ulogic;
	signal   CPMINTERCONNECTCLKEN_dly  :  std_ulogic;
	signal   CPMMCCLK_dly  :  std_ulogic;
	signal   DBGC440DEBUGHALT_dly  :  std_ulogic;
	signal   DBGC440SYSTEMSTATUS_dly  :  std_logic_vector(0 to 4);
	signal   DBGC440UNCONDDEBUGEVENT_dly  :  std_ulogic;
	signal   DCRPPCDSABUS_dly  :  std_logic_vector(0 to 9);
	signal   DCRPPCDSDBUSOUT_dly  :  std_logic_vector(0 to 31);
	signal   DCRPPCDSREAD_dly  :  std_ulogic;
	signal   DCRPPCDSWRITE_dly  :  std_ulogic;
	signal   EICC440CRITIRQ_dly  :  std_ulogic;
	signal   EICC440EXTIRQ_dly  :  std_ulogic;
	signal   FCMAPUCONFIRMINSTR_dly  :  std_ulogic;
	signal   FCMAPUCR_dly  :  std_logic_vector(0 to 3);
	signal   FCMAPUDONE_dly  :  std_ulogic;
	signal   FCMAPUEXCEPTION_dly  :  std_ulogic;
	signal   FCMAPUFPSCRFEX_dly  :  std_ulogic;
	signal   FCMAPURESULT_dly  :  std_logic_vector(0 to 31);
	signal   FCMAPURESULTVALID_dly  :  std_ulogic;
	signal   FCMAPUSLEEPNOTREADY_dly  :  std_ulogic;
	signal   FCMAPUSTOREDATA_dly  :  std_logic_vector(0 to 127);
	signal   JTGC440TCK_dly  :  std_ulogic;
	signal   JTGC440TDI_dly  :  std_ulogic;
	signal   JTGC440TMS_dly  :  std_ulogic;
	signal   JTGC440TRSTNEG_dly  :  std_ulogic;
	signal   MCMIADDRREADYTOACCEPT_dly  :  std_ulogic;
	signal   MCMIREADDATA_dly  :  std_logic_vector(0 to 127);
	signal   MCMIREADDATAERR_dly  :  std_ulogic;
	signal   MCMIREADDATAVALID_dly  :  std_ulogic;
	signal   RSTC440RESETCHIP_dly  :  std_ulogic;
	signal   RSTC440RESETCORE_dly  :  std_ulogic;
	signal   RSTC440RESETSYSTEM_dly  :  std_ulogic;
	signal   TIEC440DCURDLDCACHEPLBPRIO_dly  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDNONCACHEPLBPRIO_dly  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDTOUCHPLBPRIO_dly  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDURGENTPLBPRIO_dly  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRFLUSHPLBPRIO_dly  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRSTOREPLBPRIO_dly  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRURGENTPLBPRIO_dly  :  std_logic_vector(0 to 1);
	signal   TIEC440ENDIANRESET_dly  :  std_ulogic;
	signal   TIEC440ERPNRESET_dly  :  std_logic_vector(0 to 3);
	signal   TIEC440ICURDFETCHPLBPRIO_dly  :  std_logic_vector(0 to 1);
	signal   TIEC440ICURDSPECPLBPRIO_dly  :  std_logic_vector(0 to 1);
	signal   TIEC440ICURDTOUCHPLBPRIO_dly  :  std_logic_vector(0 to 1);
	signal   TIEC440PIR_dly  :  std_logic_vector(28 to 31);
	signal   TIEC440PVR_dly  :  std_logic_vector(28 to 31);
	signal   TIEC440USERRESET_dly  :  std_logic_vector(0 to 3);
	signal   TRCC440TRACEDISABLE_dly  :  std_ulogic;
	signal   TRCC440TRIGGEREVENTIN_dly  :  std_ulogic;

	signal   PLBPPCS0RNW_indelay  :  std_ulogic;
	signal   PLBPPCS1RNW_indelay  :  std_ulogic;
	signal   CPMDCRCLK_indelay  :  std_ulogic;
	signal   CPMDMA0LLCLK_indelay  :  std_ulogic;
	signal   CPMDMA1LLCLK_indelay  :  std_ulogic;
	signal   CPMDMA2LLCLK_indelay  :  std_ulogic;
	signal   CPMDMA3LLCLK_indelay  :  std_ulogic;
	signal   CPMINTERCONNECTCLKNTO1_indelay  :  std_ulogic;
	signal   CPMPPCMPLBCLK_indelay  :  std_ulogic;
	signal   CPMPPCS0PLBCLK_indelay  :  std_ulogic;
	signal   CPMPPCS1PLBCLK_indelay  :  std_ulogic;
	signal   DCRPPCDMACK_indelay  :  std_ulogic;
	signal   DCRPPCDMDBUSIN_indelay  :  std_logic_vector(0 to 31);
	signal   DCRPPCDMTIMEOUTWAIT_indelay  :  std_ulogic;
	signal   LLDMA0RSTENGINEREQ_indelay  :  std_ulogic;
	signal   LLDMA0RXD_indelay  :  std_logic_vector(0 to 31);
	signal   LLDMA0RXEOFN_indelay  :  std_ulogic;
	signal   LLDMA0RXEOPN_indelay  :  std_ulogic;
	signal   LLDMA0RXREM_indelay  :  std_logic_vector(0 to 3);
	signal   LLDMA0RXSOFN_indelay  :  std_ulogic;
	signal   LLDMA0RXSOPN_indelay  :  std_ulogic;
	signal   LLDMA0RXSRCRDYN_indelay  :  std_ulogic;
	signal   LLDMA0TXDSTRDYN_indelay  :  std_ulogic;
	signal   LLDMA1RSTENGINEREQ_indelay  :  std_ulogic;
	signal   LLDMA1RXD_indelay  :  std_logic_vector(0 to 31);
	signal   LLDMA1RXEOFN_indelay  :  std_ulogic;
	signal   LLDMA1RXEOPN_indelay  :  std_ulogic;
	signal   LLDMA1RXREM_indelay  :  std_logic_vector(0 to 3);
	signal   LLDMA1RXSOFN_indelay  :  std_ulogic;
	signal   LLDMA1RXSOPN_indelay  :  std_ulogic;
	signal   LLDMA1RXSRCRDYN_indelay  :  std_ulogic;
	signal   LLDMA1TXDSTRDYN_indelay  :  std_ulogic;
	signal   LLDMA2RSTENGINEREQ_indelay  :  std_ulogic;
	signal   LLDMA2RXD_indelay  :  std_logic_vector(0 to 31);
	signal   LLDMA2RXEOFN_indelay  :  std_ulogic;
	signal   LLDMA2RXEOPN_indelay  :  std_ulogic;
	signal   LLDMA2RXREM_indelay  :  std_logic_vector(0 to 3);
	signal   LLDMA2RXSOFN_indelay  :  std_ulogic;
	signal   LLDMA2RXSOPN_indelay  :  std_ulogic;
	signal   LLDMA2RXSRCRDYN_indelay  :  std_ulogic;
	signal   LLDMA2TXDSTRDYN_indelay  :  std_ulogic;
	signal   LLDMA3RSTENGINEREQ_indelay  :  std_ulogic;
	signal   LLDMA3RXD_indelay  :  std_logic_vector(0 to 31);
	signal   LLDMA3RXEOFN_indelay  :  std_ulogic;
	signal   LLDMA3RXEOPN_indelay  :  std_ulogic;
	signal   LLDMA3RXREM_indelay  :  std_logic_vector(0 to 3);
	signal   LLDMA3RXSOFN_indelay  :  std_ulogic;
	signal   LLDMA3RXSOPN_indelay  :  std_ulogic;
	signal   LLDMA3RXSRCRDYN_indelay  :  std_ulogic;
	signal   LLDMA3TXDSTRDYN_indelay  :  std_ulogic;
	signal   PLBPPCMADDRACK_indelay  :  std_ulogic;
	signal   PLBPPCMMBUSY_indelay  :  std_ulogic;
	signal   PLBPPCMMIRQ_indelay  :  std_ulogic;
	signal   PLBPPCMMRDERR_indelay  :  std_ulogic;
	signal   PLBPPCMMWRERR_indelay  :  std_ulogic;
	signal   PLBPPCMRDBTERM_indelay  :  std_ulogic;
	signal   PLBPPCMRDDACK_indelay  :  std_ulogic;
	signal   PLBPPCMRDDBUS_indelay  :  std_logic_vector(0 to 127);
	signal   PLBPPCMRDPENDPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCMRDPENDREQ_indelay  :  std_ulogic;
	signal   PLBPPCMRDWDADDR_indelay  :  std_logic_vector(0 to 3);
	signal   PLBPPCMREARBITRATE_indelay  :  std_ulogic;
	signal   PLBPPCMREQPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCMSSIZE_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCMTIMEOUT_indelay  :  std_ulogic;
	signal   PLBPPCMWRBTERM_indelay  :  std_ulogic;
	signal   PLBPPCMWRDACK_indelay  :  std_ulogic;
	signal   PLBPPCMWRPENDPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCMWRPENDREQ_indelay  :  std_ulogic;
	signal   PLBPPCS0ABORT_indelay  :  std_ulogic;
	signal   PLBPPCS0ABUS_indelay  :  std_logic_vector(0 to 31);
	signal   PLBPPCS0BE_indelay  :  std_logic_vector(0 to 15);
	signal   PLBPPCS0BUSLOCK_indelay  :  std_ulogic;
	signal   PLBPPCS0LOCKERR_indelay  :  std_ulogic;
	signal   PLBPPCS0MASTERID_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0MSIZE_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0PAVALID_indelay  :  std_ulogic;
	signal   PLBPPCS0RDBURST_indelay  :  std_ulogic;
	signal   PLBPPCS0RDPENDPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0RDPENDREQ_indelay  :  std_ulogic;
	signal   PLBPPCS0RDPRIM_indelay  :  std_ulogic;
	signal   PLBPPCS0REQPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0SAVALID_indelay  :  std_ulogic;
	signal   PLBPPCS0SIZE_indelay  :  std_logic_vector(0 to 3);
	signal   PLBPPCS0TATTRIBUTE_indelay  :  std_logic_vector(0 to 15);
	signal   PLBPPCS0TYPE_indelay  :  std_logic_vector(0 to 2);
	signal   PLBPPCS0UABUS_indelay  :  std_logic_vector(28 to 31);
	signal   PLBPPCS0WRBURST_indelay  :  std_ulogic;
	signal   PLBPPCS0WRDBUS_indelay  :  std_logic_vector(0 to 127);
	signal   PLBPPCS0WRPENDPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS0WRPENDREQ_indelay  :  std_ulogic;
	signal   PLBPPCS0WRPRIM_indelay  :  std_ulogic;
	signal   PLBPPCS1ABORT_indelay  :  std_ulogic;
	signal   PLBPPCS1ABUS_indelay  :  std_logic_vector(0 to 31);
	signal   PLBPPCS1BE_indelay  :  std_logic_vector(0 to 15);
	signal   PLBPPCS1BUSLOCK_indelay  :  std_ulogic;
	signal   PLBPPCS1LOCKERR_indelay  :  std_ulogic;
	signal   PLBPPCS1MASTERID_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1MSIZE_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1PAVALID_indelay  :  std_ulogic;
	signal   PLBPPCS1RDBURST_indelay  :  std_ulogic;
	signal   PLBPPCS1RDPENDPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1RDPENDREQ_indelay  :  std_ulogic;
	signal   PLBPPCS1RDPRIM_indelay  :  std_ulogic;
	signal   PLBPPCS1REQPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1SAVALID_indelay  :  std_ulogic;
	signal   PLBPPCS1SIZE_indelay  :  std_logic_vector(0 to 3);
	signal   PLBPPCS1TATTRIBUTE_indelay  :  std_logic_vector(0 to 15);
	signal   PLBPPCS1TYPE_indelay  :  std_logic_vector(0 to 2);
	signal   PLBPPCS1UABUS_indelay  :  std_logic_vector(28 to 31);
	signal   PLBPPCS1WRBURST_indelay  :  std_ulogic;
	signal   PLBPPCS1WRDBUS_indelay  :  std_logic_vector(0 to 127);
	signal   PLBPPCS1WRPENDPRI_indelay  :  std_logic_vector(0 to 1);
	signal   PLBPPCS1WRPENDREQ_indelay  :  std_ulogic;
	signal   PLBPPCS1WRPRIM_indelay  :  std_ulogic;
	signal   TIEDCRBASEADDR_indelay  :  std_logic_vector(0 to 1);
	signal   CPMC440CLK_indelay  :  std_ulogic;
	signal   CPMC440CLKEN_indelay  :  std_ulogic;
	signal   CPMC440CORECLOCKINACTIVE_indelay  :  std_ulogic;
	signal   CPMC440TIMERCLOCK_indelay  :  std_ulogic;
	signal   CPMFCMCLK_indelay  :  std_ulogic;
	signal   CPMINTERCONNECTCLK_indelay  :  std_ulogic;
	signal   CPMINTERCONNECTCLKEN_indelay  :  std_ulogic;
	signal   CPMMCCLK_indelay  :  std_ulogic;
	signal   DBGC440DEBUGHALT_indelay  :  std_ulogic;
	signal   DBGC440SYSTEMSTATUS_indelay  :  std_logic_vector(0 to 4);
	signal   DBGC440UNCONDDEBUGEVENT_indelay  :  std_ulogic;
	signal   DCRPPCDSABUS_indelay  :  std_logic_vector(0 to 9);
	signal   DCRPPCDSDBUSOUT_indelay  :  std_logic_vector(0 to 31);
	signal   DCRPPCDSREAD_indelay  :  std_ulogic;
	signal   DCRPPCDSWRITE_indelay  :  std_ulogic;
	signal   EICC440CRITIRQ_indelay  :  std_ulogic;
	signal   EICC440EXTIRQ_indelay  :  std_ulogic;
	signal   FCMAPUCONFIRMINSTR_indelay  :  std_ulogic;
	signal   FCMAPUCR_indelay  :  std_logic_vector(0 to 3);
	signal   FCMAPUDONE_indelay  :  std_ulogic;
	signal   FCMAPUEXCEPTION_indelay  :  std_ulogic;
	signal   FCMAPUFPSCRFEX_indelay  :  std_ulogic;
	signal   FCMAPURESULT_indelay  :  std_logic_vector(0 to 31);
	signal   FCMAPURESULTVALID_indelay  :  std_ulogic;
	signal   FCMAPUSLEEPNOTREADY_indelay  :  std_ulogic;
	signal   FCMAPUSTOREDATA_indelay  :  std_logic_vector(0 to 127);
	signal   JTGC440TCK_indelay  :  std_ulogic;
	signal   JTGC440TDI_indelay  :  std_ulogic;
	signal   JTGC440TMS_indelay  :  std_ulogic;
	signal   JTGC440TRSTNEG_indelay  :  std_ulogic;
	signal   MCMIADDRREADYTOACCEPT_indelay  :  std_ulogic;
	signal   MCMIREADDATA_indelay  :  std_logic_vector(0 to 127);
	signal   MCMIREADDATAERR_indelay  :  std_ulogic;
	signal   MCMIREADDATAVALID_indelay  :  std_ulogic;
	signal   RSTC440RESETCHIP_indelay  :  std_ulogic;
	signal   RSTC440RESETCORE_indelay  :  std_ulogic;
	signal   RSTC440RESETSYSTEM_indelay  :  std_ulogic;
	signal   TIEC440DCURDLDCACHEPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDNONCACHEPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDTOUCHPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440DCURDURGENTPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRFLUSHPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRSTOREPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440DCUWRURGENTPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440ENDIANRESET_indelay  :  std_ulogic;
	signal   TIEC440ERPNRESET_indelay  :  std_logic_vector(0 to 3);
	signal   TIEC440ICURDFETCHPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440ICURDSPECPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440ICURDTOUCHPLBPRIO_indelay  :  std_logic_vector(0 to 1);
	signal   TIEC440PIR_indelay  :  std_logic_vector(28 to 31);
	signal   TIEC440PVR_indelay  :  std_logic_vector(28 to 31);
	signal   TIEC440USERRESET_indelay  :  std_logic_vector(0 to 3);
	signal   TRCC440TRACEDISABLE_indelay  :  std_ulogic;
	signal   TRCC440TRIGGEREVENTIN_indelay  :  std_ulogic;

begin
	WireDelay : block
	begin
              VitalWireDelay (PLBPPCS0RNW_ipd,PLBPPCS0RNW,tipd_PLBPPCS0RNW);
              VitalWireDelay (PLBPPCS1RNW_ipd,PLBPPCS1RNW,tipd_PLBPPCS1RNW);
              VitalWireDelay (CPMDCRCLK_ipd,CPMDCRCLK,tipd_CPMDCRCLK);
              VitalWireDelay (CPMDMA0LLCLK_ipd,CPMDMA0LLCLK,tipd_CPMDMA0LLCLK);
              VitalWireDelay (CPMDMA1LLCLK_ipd,CPMDMA1LLCLK,tipd_CPMDMA1LLCLK);
              VitalWireDelay (CPMDMA2LLCLK_ipd,CPMDMA2LLCLK,tipd_CPMDMA2LLCLK);
              VitalWireDelay (CPMDMA3LLCLK_ipd,CPMDMA3LLCLK,tipd_CPMDMA3LLCLK);
              VitalWireDelay (CPMINTERCONNECTCLKNTO1_ipd,CPMINTERCONNECTCLKNTO1,tipd_CPMINTERCONNECTCLKNTO1);
              VitalWireDelay (CPMPPCMPLBCLK_ipd,CPMPPCMPLBCLK,tipd_CPMPPCMPLBCLK);
              VitalWireDelay (CPMPPCS0PLBCLK_ipd,CPMPPCS0PLBCLK,tipd_CPMPPCS0PLBCLK);
              VitalWireDelay (CPMPPCS1PLBCLK_ipd,CPMPPCS1PLBCLK,tipd_CPMPPCS1PLBCLK);
              VitalWireDelay (DCRPPCDMACK_ipd,DCRPPCDMACK,tipd_DCRPPCDMACK);
           DCRPPCDMDBUSIN_DELAY : for i in 0 to 31 generate
              VitalWireDelay (DCRPPCDMDBUSIN_ipd(i),DCRPPCDMDBUSIN(i),tipd_DCRPPCDMDBUSIN(i));
           end generate DCRPPCDMDBUSIN_DELAY;
              VitalWireDelay (DCRPPCDMTIMEOUTWAIT_ipd,DCRPPCDMTIMEOUTWAIT,tipd_DCRPPCDMTIMEOUTWAIT);
              VitalWireDelay (LLDMA0RSTENGINEREQ_ipd,LLDMA0RSTENGINEREQ,tipd_LLDMA0RSTENGINEREQ);
           LLDMA0RXD_DELAY : for i in 0 to 31 generate
              VitalWireDelay (LLDMA0RXD_ipd(i),LLDMA0RXD(i),tipd_LLDMA0RXD(i));
           end generate LLDMA0RXD_DELAY;
              VitalWireDelay (LLDMA0RXEOFN_ipd,LLDMA0RXEOFN,tipd_LLDMA0RXEOFN);
              VitalWireDelay (LLDMA0RXEOPN_ipd,LLDMA0RXEOPN,tipd_LLDMA0RXEOPN);
           LLDMA0RXREM_DELAY : for i in 0 to 3 generate
              VitalWireDelay (LLDMA0RXREM_ipd(i),LLDMA0RXREM(i),tipd_LLDMA0RXREM(i));
           end generate LLDMA0RXREM_DELAY;
              VitalWireDelay (LLDMA0RXSOFN_ipd,LLDMA0RXSOFN,tipd_LLDMA0RXSOFN);
              VitalWireDelay (LLDMA0RXSOPN_ipd,LLDMA0RXSOPN,tipd_LLDMA0RXSOPN);
              VitalWireDelay (LLDMA0RXSRCRDYN_ipd,LLDMA0RXSRCRDYN,tipd_LLDMA0RXSRCRDYN);
              VitalWireDelay (LLDMA0TXDSTRDYN_ipd,LLDMA0TXDSTRDYN,tipd_LLDMA0TXDSTRDYN);
              VitalWireDelay (LLDMA1RSTENGINEREQ_ipd,LLDMA1RSTENGINEREQ,tipd_LLDMA1RSTENGINEREQ);
           LLDMA1RXD_DELAY : for i in 0 to 31 generate
              VitalWireDelay (LLDMA1RXD_ipd(i),LLDMA1RXD(i),tipd_LLDMA1RXD(i));
           end generate LLDMA1RXD_DELAY;
              VitalWireDelay (LLDMA1RXEOFN_ipd,LLDMA1RXEOFN,tipd_LLDMA1RXEOFN);
              VitalWireDelay (LLDMA1RXEOPN_ipd,LLDMA1RXEOPN,tipd_LLDMA1RXEOPN);
           LLDMA1RXREM_DELAY : for i in 0 to 3 generate
              VitalWireDelay (LLDMA1RXREM_ipd(i),LLDMA1RXREM(i),tipd_LLDMA1RXREM(i));
           end generate LLDMA1RXREM_DELAY;
              VitalWireDelay (LLDMA1RXSOFN_ipd,LLDMA1RXSOFN,tipd_LLDMA1RXSOFN);
              VitalWireDelay (LLDMA1RXSOPN_ipd,LLDMA1RXSOPN,tipd_LLDMA1RXSOPN);
              VitalWireDelay (LLDMA1RXSRCRDYN_ipd,LLDMA1RXSRCRDYN,tipd_LLDMA1RXSRCRDYN);
              VitalWireDelay (LLDMA1TXDSTRDYN_ipd,LLDMA1TXDSTRDYN,tipd_LLDMA1TXDSTRDYN);
              VitalWireDelay (LLDMA2RSTENGINEREQ_ipd,LLDMA2RSTENGINEREQ,tipd_LLDMA2RSTENGINEREQ);
           LLDMA2RXD_DELAY : for i in 0 to 31 generate
              VitalWireDelay (LLDMA2RXD_ipd(i),LLDMA2RXD(i),tipd_LLDMA2RXD(i));
           end generate LLDMA2RXD_DELAY;
              VitalWireDelay (LLDMA2RXEOFN_ipd,LLDMA2RXEOFN,tipd_LLDMA2RXEOFN);
              VitalWireDelay (LLDMA2RXEOPN_ipd,LLDMA2RXEOPN,tipd_LLDMA2RXEOPN);
           LLDMA2RXREM_DELAY : for i in 0 to 3 generate
              VitalWireDelay (LLDMA2RXREM_ipd(i),LLDMA2RXREM(i),tipd_LLDMA2RXREM(i));
           end generate LLDMA2RXREM_DELAY;
              VitalWireDelay (LLDMA2RXSOFN_ipd,LLDMA2RXSOFN,tipd_LLDMA2RXSOFN);
              VitalWireDelay (LLDMA2RXSOPN_ipd,LLDMA2RXSOPN,tipd_LLDMA2RXSOPN);
              VitalWireDelay (LLDMA2RXSRCRDYN_ipd,LLDMA2RXSRCRDYN,tipd_LLDMA2RXSRCRDYN);
              VitalWireDelay (LLDMA2TXDSTRDYN_ipd,LLDMA2TXDSTRDYN,tipd_LLDMA2TXDSTRDYN);
              VitalWireDelay (LLDMA3RSTENGINEREQ_ipd,LLDMA3RSTENGINEREQ,tipd_LLDMA3RSTENGINEREQ);
           LLDMA3RXD_DELAY : for i in 0 to 31 generate
              VitalWireDelay (LLDMA3RXD_ipd(i),LLDMA3RXD(i),tipd_LLDMA3RXD(i));
           end generate LLDMA3RXD_DELAY;
              VitalWireDelay (LLDMA3RXEOFN_ipd,LLDMA3RXEOFN,tipd_LLDMA3RXEOFN);
              VitalWireDelay (LLDMA3RXEOPN_ipd,LLDMA3RXEOPN,tipd_LLDMA3RXEOPN);
           LLDMA3RXREM_DELAY : for i in 0 to 3 generate
              VitalWireDelay (LLDMA3RXREM_ipd(i),LLDMA3RXREM(i),tipd_LLDMA3RXREM(i));
           end generate LLDMA3RXREM_DELAY;
              VitalWireDelay (LLDMA3RXSOFN_ipd,LLDMA3RXSOFN,tipd_LLDMA3RXSOFN);
              VitalWireDelay (LLDMA3RXSOPN_ipd,LLDMA3RXSOPN,tipd_LLDMA3RXSOPN);
              VitalWireDelay (LLDMA3RXSRCRDYN_ipd,LLDMA3RXSRCRDYN,tipd_LLDMA3RXSRCRDYN);
              VitalWireDelay (LLDMA3TXDSTRDYN_ipd,LLDMA3TXDSTRDYN,tipd_LLDMA3TXDSTRDYN);
              VitalWireDelay (PLBPPCMADDRACK_ipd,PLBPPCMADDRACK,tipd_PLBPPCMADDRACK);
              VitalWireDelay (PLBPPCMMBUSY_ipd,PLBPPCMMBUSY,tipd_PLBPPCMMBUSY);
              VitalWireDelay (PLBPPCMMIRQ_ipd,PLBPPCMMIRQ,tipd_PLBPPCMMIRQ);
              VitalWireDelay (PLBPPCMMRDERR_ipd,PLBPPCMMRDERR,tipd_PLBPPCMMRDERR);
              VitalWireDelay (PLBPPCMMWRERR_ipd,PLBPPCMMWRERR,tipd_PLBPPCMMWRERR);
              VitalWireDelay (PLBPPCMRDBTERM_ipd,PLBPPCMRDBTERM,tipd_PLBPPCMRDBTERM);
              VitalWireDelay (PLBPPCMRDDACK_ipd,PLBPPCMRDDACK,tipd_PLBPPCMRDDACK);
           PLBPPCMRDDBUS_DELAY : for i in 0 to 127 generate
              VitalWireDelay (PLBPPCMRDDBUS_ipd(i),PLBPPCMRDDBUS(i),tipd_PLBPPCMRDDBUS(i));
           end generate PLBPPCMRDDBUS_DELAY;
           PLBPPCMRDPENDPRI_DELAY : for i in 0 to 1 generate
              VitalWireDelay (PLBPPCMRDPENDPRI_ipd(i),PLBPPCMRDPENDPRI(i),tipd_PLBPPCMRDPENDPRI(i));
           end generate PLBPPCMRDPENDPRI_DELAY;
              VitalWireDelay (PLBPPCMRDPENDREQ_ipd,PLBPPCMRDPENDREQ,tipd_PLBPPCMRDPENDREQ);
           PLBPPCMRDWDADDR_DELAY : for i in 0 to 3 generate
              VitalWireDelay (PLBPPCMRDWDADDR_ipd(i),PLBPPCMRDWDADDR(i),tipd_PLBPPCMRDWDADDR(i));
           end generate PLBPPCMRDWDADDR_DELAY;
              VitalWireDelay (PLBPPCMREARBITRATE_ipd,PLBPPCMREARBITRATE,tipd_PLBPPCMREARBITRATE);
           PLBPPCMREQPRI_DELAY : for i in 0 to 1 generate
              VitalWireDelay (PLBPPCMREQPRI_ipd(i),PLBPPCMREQPRI(i),tipd_PLBPPCMREQPRI(i));
           end generate PLBPPCMREQPRI_DELAY;
           PLBPPCMSSIZE_DELAY : for i in 0 to 1 generate
              VitalWireDelay (PLBPPCMSSIZE_ipd(i),PLBPPCMSSIZE(i),tipd_PLBPPCMSSIZE(i));
           end generate PLBPPCMSSIZE_DELAY;
              VitalWireDelay (PLBPPCMTIMEOUT_ipd,PLBPPCMTIMEOUT,tipd_PLBPPCMTIMEOUT);
              VitalWireDelay (PLBPPCMWRBTERM_ipd,PLBPPCMWRBTERM,tipd_PLBPPCMWRBTERM);
              VitalWireDelay (PLBPPCMWRDACK_ipd,PLBPPCMWRDACK,tipd_PLBPPCMWRDACK);
           PLBPPCMWRPENDPRI_DELAY : for i in 0 to 1 generate
              VitalWireDelay (PLBPPCMWRPENDPRI_ipd(i),PLBPPCMWRPENDPRI(i),tipd_PLBPPCMWRPENDPRI(i));
           end generate PLBPPCMWRPENDPRI_DELAY;
              VitalWireDelay (PLBPPCMWRPENDREQ_ipd,PLBPPCMWRPENDREQ,tipd_PLBPPCMWRPENDREQ);
              VitalWireDelay (PLBPPCS0ABORT_ipd,PLBPPCS0ABORT,tipd_PLBPPCS0ABORT);
           PLBPPCS0ABUS_DELAY : for i in 0 to 31 generate
              VitalWireDelay (PLBPPCS0ABUS_ipd(i),PLBPPCS0ABUS(i),tipd_PLBPPCS0ABUS(i));
           end generate PLBPPCS0ABUS_DELAY;
           PLBPPCS0BE_DELAY : for i in 0 to 15 generate
              VitalWireDelay (PLBPPCS0BE_ipd(i),PLBPPCS0BE(i),tipd_PLBPPCS0BE(i));
           end generate PLBPPCS0BE_DELAY;
              VitalWireDelay (PLBPPCS0BUSLOCK_ipd,PLBPPCS0BUSLOCK,tipd_PLBPPCS0BUSLOCK);
              VitalWireDelay (PLBPPCS0LOCKERR_ipd,PLBPPCS0LOCKERR,tipd_PLBPPCS0LOCKERR);
           PLBPPCS0MASTERID_DELAY : for i in 0 to 1 generate
              VitalWireDelay (PLBPPCS0MASTERID_ipd(i),PLBPPCS0MASTERID(i),tipd_PLBPPCS0MASTERID(i));
           end generate PLBPPCS0MASTERID_DELAY;
           PLBPPCS0MSIZE_DELAY : for i in 0 to 1 generate
              VitalWireDelay (PLBPPCS0MSIZE_ipd(i),PLBPPCS0MSIZE(i),tipd_PLBPPCS0MSIZE(i));
           end generate PLBPPCS0MSIZE_DELAY;
              VitalWireDelay (PLBPPCS0PAVALID_ipd,PLBPPCS0PAVALID,tipd_PLBPPCS0PAVALID);
              VitalWireDelay (PLBPPCS0RDBURST_ipd,PLBPPCS0RDBURST,tipd_PLBPPCS0RDBURST);
           PLBPPCS0RDPENDPRI_DELAY : for i in 0 to 1 generate
              VitalWireDelay (PLBPPCS0RDPENDPRI_ipd(i),PLBPPCS0RDPENDPRI(i),tipd_PLBPPCS0RDPENDPRI(i));
           end generate PLBPPCS0RDPENDPRI_DELAY;
              VitalWireDelay (PLBPPCS0RDPENDREQ_ipd,PLBPPCS0RDPENDREQ,tipd_PLBPPCS0RDPENDREQ);
              VitalWireDelay (PLBPPCS0RDPRIM_ipd,PLBPPCS0RDPRIM,tipd_PLBPPCS0RDPRIM);
           PLBPPCS0REQPRI_DELAY : for i in 0 to 1 generate
              VitalWireDelay (PLBPPCS0REQPRI_ipd(i),PLBPPCS0REQPRI(i),tipd_PLBPPCS0REQPRI(i));
           end generate PLBPPCS0REQPRI_DELAY;
              VitalWireDelay (PLBPPCS0SAVALID_ipd,PLBPPCS0SAVALID,tipd_PLBPPCS0SAVALID);
           PLBPPCS0SIZE_DELAY : for i in 0 to 3 generate
              VitalWireDelay (PLBPPCS0SIZE_ipd(i),PLBPPCS0SIZE(i),tipd_PLBPPCS0SIZE(i));
           end generate PLBPPCS0SIZE_DELAY;
           PLBPPCS0TATTRIBUTE_DELAY : for i in 0 to 15 generate
              VitalWireDelay (PLBPPCS0TATTRIBUTE_ipd(i),PLBPPCS0TATTRIBUTE(i),tipd_PLBPPCS0TATTRIBUTE(i));
           end generate PLBPPCS0TATTRIBUTE_DELAY;
           PLBPPCS0TYPE_DELAY : for i in 0 to 2 generate
              VitalWireDelay (PLBPPCS0TYPE_ipd(i),PLBPPCS0TYPE(i),tipd_PLBPPCS0TYPE(i));
           end generate PLBPPCS0TYPE_DELAY;
           PLBPPCS0UABUS_DELAY : for i in 28 to 31 generate
              VitalWireDelay (PLBPPCS0UABUS_ipd(i),PLBPPCS0UABUS(i),tipd_PLBPPCS0UABUS(i));
           end generate PLBPPCS0UABUS_DELAY;
              VitalWireDelay (PLBPPCS0WRBURST_ipd,PLBPPCS0WRBURST,tipd_PLBPPCS0WRBURST);
           PLBPPCS0WRDBUS_DELAY : for i in 0 to 127 generate
              VitalWireDelay (PLBPPCS0WRDBUS_ipd(i),PLBPPCS0WRDBUS(i),tipd_PLBPPCS0WRDBUS(i));
           end generate PLBPPCS0WRDBUS_DELAY;
           PLBPPCS0WRPENDPRI_DELAY : for i in 0 to 1 generate
              VitalWireDelay (PLBPPCS0WRPENDPRI_ipd(i),PLBPPCS0WRPENDPRI(i),tipd_PLBPPCS0WRPENDPRI(i));
           end generate PLBPPCS0WRPENDPRI_DELAY;
              VitalWireDelay (PLBPPCS0WRPENDREQ_ipd,PLBPPCS0WRPENDREQ,tipd_PLBPPCS0WRPENDREQ);
              VitalWireDelay (PLBPPCS0WRPRIM_ipd,PLBPPCS0WRPRIM,tipd_PLBPPCS0WRPRIM);
              VitalWireDelay (PLBPPCS1ABORT_ipd,PLBPPCS1ABORT,tipd_PLBPPCS1ABORT);
           PLBPPCS1ABUS_DELAY : for i in 0 to 31 generate
              VitalWireDelay (PLBPPCS1ABUS_ipd(i),PLBPPCS1ABUS(i),tipd_PLBPPCS1ABUS(i));
           end generate PLBPPCS1ABUS_DELAY;
           PLBPPCS1BE_DELAY : for i in 0 to 15 generate
              VitalWireDelay (PLBPPCS1BE_ipd(i),PLBPPCS1BE(i),tipd_PLBPPCS1BE(i));
           end generate PLBPPCS1BE_DELAY;
              VitalWireDelay (PLBPPCS1BUSLOCK_ipd,PLBPPCS1BUSLOCK,tipd_PLBPPCS1BUSLOCK);
              VitalWireDelay (PLBPPCS1LOCKERR_ipd,PLBPPCS1LOCKERR,tipd_PLBPPCS1LOCKERR);
           PLBPPCS1MASTERID_DELAY : for i in 0 to 1 generate
              VitalWireDelay (PLBPPCS1MASTERID_ipd(i),PLBPPCS1MASTERID(i),tipd_PLBPPCS1MASTERID(i));
           end generate PLBPPCS1MASTERID_DELAY;
           PLBPPCS1MSIZE_DELAY : for i in 0 to 1 generate
              VitalWireDelay (PLBPPCS1MSIZE_ipd(i),PLBPPCS1MSIZE(i),tipd_PLBPPCS1MSIZE(i));
           end generate PLBPPCS1MSIZE_DELAY;
              VitalWireDelay (PLBPPCS1PAVALID_ipd,PLBPPCS1PAVALID,tipd_PLBPPCS1PAVALID);
              VitalWireDelay (PLBPPCS1RDBURST_ipd,PLBPPCS1RDBURST,tipd_PLBPPCS1RDBURST);
           PLBPPCS1RDPENDPRI_DELAY : for i in 0 to 1 generate
              VitalWireDelay (PLBPPCS1RDPENDPRI_ipd(i),PLBPPCS1RDPENDPRI(i),tipd_PLBPPCS1RDPENDPRI(i));
           end generate PLBPPCS1RDPENDPRI_DELAY;
              VitalWireDelay (PLBPPCS1RDPENDREQ_ipd,PLBPPCS1RDPENDREQ,tipd_PLBPPCS1RDPENDREQ);
              VitalWireDelay (PLBPPCS1RDPRIM_ipd,PLBPPCS1RDPRIM,tipd_PLBPPCS1RDPRIM);
           PLBPPCS1REQPRI_DELAY : for i in 0 to 1 generate
              VitalWireDelay (PLBPPCS1REQPRI_ipd(i),PLBPPCS1REQPRI(i),tipd_PLBPPCS1REQPRI(i));
           end generate PLBPPCS1REQPRI_DELAY;
              VitalWireDelay (PLBPPCS1SAVALID_ipd,PLBPPCS1SAVALID,tipd_PLBPPCS1SAVALID);
           PLBPPCS1SIZE_DELAY : for i in 0 to 3 generate
              VitalWireDelay (PLBPPCS1SIZE_ipd(i),PLBPPCS1SIZE(i),tipd_PLBPPCS1SIZE(i));
           end generate PLBPPCS1SIZE_DELAY;
           PLBPPCS1TATTRIBUTE_DELAY : for i in 0 to 15 generate
              VitalWireDelay (PLBPPCS1TATTRIBUTE_ipd(i),PLBPPCS1TATTRIBUTE(i),tipd_PLBPPCS1TATTRIBUTE(i));
           end generate PLBPPCS1TATTRIBUTE_DELAY;
           PLBPPCS1TYPE_DELAY : for i in 0 to 2 generate
              VitalWireDelay (PLBPPCS1TYPE_ipd(i),PLBPPCS1TYPE(i),tipd_PLBPPCS1TYPE(i));
           end generate PLBPPCS1TYPE_DELAY;
           PLBPPCS1UABUS_DELAY : for i in 28 to 31 generate
              VitalWireDelay (PLBPPCS1UABUS_ipd(i),PLBPPCS1UABUS(i),tipd_PLBPPCS1UABUS(i));
           end generate PLBPPCS1UABUS_DELAY;
              VitalWireDelay (PLBPPCS1WRBURST_ipd,PLBPPCS1WRBURST,tipd_PLBPPCS1WRBURST);
           PLBPPCS1WRDBUS_DELAY : for i in 0 to 127 generate
              VitalWireDelay (PLBPPCS1WRDBUS_ipd(i),PLBPPCS1WRDBUS(i),tipd_PLBPPCS1WRDBUS(i));
           end generate PLBPPCS1WRDBUS_DELAY;
           PLBPPCS1WRPENDPRI_DELAY : for i in 0 to 1 generate
              VitalWireDelay (PLBPPCS1WRPENDPRI_ipd(i),PLBPPCS1WRPENDPRI(i),tipd_PLBPPCS1WRPENDPRI(i));
           end generate PLBPPCS1WRPENDPRI_DELAY;
              VitalWireDelay (PLBPPCS1WRPENDREQ_ipd,PLBPPCS1WRPENDREQ,tipd_PLBPPCS1WRPENDREQ);
              VitalWireDelay (PLBPPCS1WRPRIM_ipd,PLBPPCS1WRPRIM,tipd_PLBPPCS1WRPRIM);
           TIEDCRBASEADDR_DELAY : for i in 0 to 1 generate
              VitalWireDelay (TIEDCRBASEADDR_ipd(i),TIEDCRBASEADDR(i),tipd_TIEDCRBASEADDR(i));
           end generate TIEDCRBASEADDR_DELAY;
              VitalWireDelay (CPMC440CLK_ipd,CPMC440CLK,tipd_CPMC440CLK);
              VitalWireDelay (CPMC440CLKEN_ipd,CPMC440CLKEN,tipd_CPMC440CLKEN);
              VitalWireDelay (CPMC440CORECLOCKINACTIVE_ipd,CPMC440CORECLOCKINACTIVE,tipd_CPMC440CORECLOCKINACTIVE);
              VitalWireDelay (CPMC440TIMERCLOCK_ipd,CPMC440TIMERCLOCK,tipd_CPMC440TIMERCLOCK);
              VitalWireDelay (CPMFCMCLK_ipd,CPMFCMCLK,tipd_CPMFCMCLK);
              VitalWireDelay (CPMINTERCONNECTCLK_ipd,CPMINTERCONNECTCLK,tipd_CPMINTERCONNECTCLK);
              VitalWireDelay (CPMINTERCONNECTCLKEN_ipd,CPMINTERCONNECTCLKEN,tipd_CPMINTERCONNECTCLKEN);
              VitalWireDelay (CPMMCCLK_ipd,CPMMCCLK,tipd_CPMMCCLK);
              VitalWireDelay (DBGC440DEBUGHALT_ipd,DBGC440DEBUGHALT,tipd_DBGC440DEBUGHALT);
           DBGC440SYSTEMSTATUS_DELAY : for i in 0 to 4 generate
              VitalWireDelay (DBGC440SYSTEMSTATUS_ipd(i),DBGC440SYSTEMSTATUS(i),tipd_DBGC440SYSTEMSTATUS(i));
           end generate DBGC440SYSTEMSTATUS_DELAY;
              VitalWireDelay (DBGC440UNCONDDEBUGEVENT_ipd,DBGC440UNCONDDEBUGEVENT,tipd_DBGC440UNCONDDEBUGEVENT);
           DCRPPCDSABUS_DELAY : for i in 0 to 9 generate
              VitalWireDelay (DCRPPCDSABUS_ipd(i),DCRPPCDSABUS(i),tipd_DCRPPCDSABUS(i));
           end generate DCRPPCDSABUS_DELAY;
           DCRPPCDSDBUSOUT_DELAY : for i in 0 to 31 generate
              VitalWireDelay (DCRPPCDSDBUSOUT_ipd(i),DCRPPCDSDBUSOUT(i),tipd_DCRPPCDSDBUSOUT(i));
           end generate DCRPPCDSDBUSOUT_DELAY;
              VitalWireDelay (DCRPPCDSREAD_ipd,DCRPPCDSREAD,tipd_DCRPPCDSREAD);
              VitalWireDelay (DCRPPCDSWRITE_ipd,DCRPPCDSWRITE,tipd_DCRPPCDSWRITE);
              VitalWireDelay (EICC440CRITIRQ_ipd,EICC440CRITIRQ,tipd_EICC440CRITIRQ);
              VitalWireDelay (EICC440EXTIRQ_ipd,EICC440EXTIRQ,tipd_EICC440EXTIRQ);
              VitalWireDelay (FCMAPUCONFIRMINSTR_ipd,FCMAPUCONFIRMINSTR,tipd_FCMAPUCONFIRMINSTR);
           FCMAPUCR_DELAY : for i in 0 to 3 generate
              VitalWireDelay (FCMAPUCR_ipd(i),FCMAPUCR(i),tipd_FCMAPUCR(i));
           end generate FCMAPUCR_DELAY;
              VitalWireDelay (FCMAPUDONE_ipd,FCMAPUDONE,tipd_FCMAPUDONE);
              VitalWireDelay (FCMAPUEXCEPTION_ipd,FCMAPUEXCEPTION,tipd_FCMAPUEXCEPTION);
              VitalWireDelay (FCMAPUFPSCRFEX_ipd,FCMAPUFPSCRFEX,tipd_FCMAPUFPSCRFEX);
           FCMAPURESULT_DELAY : for i in 0 to 31 generate
              VitalWireDelay (FCMAPURESULT_ipd(i),FCMAPURESULT(i),tipd_FCMAPURESULT(i));
           end generate FCMAPURESULT_DELAY;
              VitalWireDelay (FCMAPURESULTVALID_ipd,FCMAPURESULTVALID,tipd_FCMAPURESULTVALID);
              VitalWireDelay (FCMAPUSLEEPNOTREADY_ipd,FCMAPUSLEEPNOTREADY,tipd_FCMAPUSLEEPNOTREADY);
           FCMAPUSTOREDATA_DELAY : for i in 0 to 127 generate
              VitalWireDelay (FCMAPUSTOREDATA_ipd(i),FCMAPUSTOREDATA(i),tipd_FCMAPUSTOREDATA(i));
           end generate FCMAPUSTOREDATA_DELAY;
              VitalWireDelay (JTGC440TCK_ipd,JTGC440TCK,tipd_JTGC440TCK);
              VitalWireDelay (JTGC440TDI_ipd,JTGC440TDI,tipd_JTGC440TDI);
              VitalWireDelay (JTGC440TMS_ipd,JTGC440TMS,tipd_JTGC440TMS);
              VitalWireDelay (JTGC440TRSTNEG_ipd,JTGC440TRSTNEG,tipd_JTGC440TRSTNEG);
              VitalWireDelay (MCMIADDRREADYTOACCEPT_ipd,MCMIADDRREADYTOACCEPT,tipd_MCMIADDRREADYTOACCEPT);
           MCMIREADDATA_DELAY : for i in 0 to 127 generate
              VitalWireDelay (MCMIREADDATA_ipd(i),MCMIREADDATA(i),tipd_MCMIREADDATA(i));
           end generate MCMIREADDATA_DELAY;
              VitalWireDelay (MCMIREADDATAERR_ipd,MCMIREADDATAERR,tipd_MCMIREADDATAERR);
              VitalWireDelay (MCMIREADDATAVALID_ipd,MCMIREADDATAVALID,tipd_MCMIREADDATAVALID);
              VitalWireDelay (RSTC440RESETCHIP_ipd,RSTC440RESETCHIP,tipd_RSTC440RESETCHIP);
              VitalWireDelay (RSTC440RESETCORE_ipd,RSTC440RESETCORE,tipd_RSTC440RESETCORE);
              VitalWireDelay (RSTC440RESETSYSTEM_ipd,RSTC440RESETSYSTEM,tipd_RSTC440RESETSYSTEM);
           TIEC440DCURDLDCACHEPLBPRIO_DELAY : for i in 0 to 1 generate
              VitalWireDelay (TIEC440DCURDLDCACHEPLBPRIO_ipd(i),TIEC440DCURDLDCACHEPLBPRIO(i),tipd_TIEC440DCURDLDCACHEPLBPRIO(i));
           end generate TIEC440DCURDLDCACHEPLBPRIO_DELAY;
           TIEC440DCURDNONCACHEPLBPRIO_DELAY : for i in 0 to 1 generate
              VitalWireDelay (TIEC440DCURDNONCACHEPLBPRIO_ipd(i),TIEC440DCURDNONCACHEPLBPRIO(i),tipd_TIEC440DCURDNONCACHEPLBPRIO(i));
           end generate TIEC440DCURDNONCACHEPLBPRIO_DELAY;
           TIEC440DCURDTOUCHPLBPRIO_DELAY : for i in 0 to 1 generate
              VitalWireDelay (TIEC440DCURDTOUCHPLBPRIO_ipd(i),TIEC440DCURDTOUCHPLBPRIO(i),tipd_TIEC440DCURDTOUCHPLBPRIO(i));
           end generate TIEC440DCURDTOUCHPLBPRIO_DELAY;
           TIEC440DCURDURGENTPLBPRIO_DELAY : for i in 0 to 1 generate
              VitalWireDelay (TIEC440DCURDURGENTPLBPRIO_ipd(i),TIEC440DCURDURGENTPLBPRIO(i),tipd_TIEC440DCURDURGENTPLBPRIO(i));
           end generate TIEC440DCURDURGENTPLBPRIO_DELAY;
           TIEC440DCUWRFLUSHPLBPRIO_DELAY : for i in 0 to 1 generate
              VitalWireDelay (TIEC440DCUWRFLUSHPLBPRIO_ipd(i),TIEC440DCUWRFLUSHPLBPRIO(i),tipd_TIEC440DCUWRFLUSHPLBPRIO(i));
           end generate TIEC440DCUWRFLUSHPLBPRIO_DELAY;
           TIEC440DCUWRSTOREPLBPRIO_DELAY : for i in 0 to 1 generate
              VitalWireDelay (TIEC440DCUWRSTOREPLBPRIO_ipd(i),TIEC440DCUWRSTOREPLBPRIO(i),tipd_TIEC440DCUWRSTOREPLBPRIO(i));
           end generate TIEC440DCUWRSTOREPLBPRIO_DELAY;
           TIEC440DCUWRURGENTPLBPRIO_DELAY : for i in 0 to 1 generate
              VitalWireDelay (TIEC440DCUWRURGENTPLBPRIO_ipd(i),TIEC440DCUWRURGENTPLBPRIO(i),tipd_TIEC440DCUWRURGENTPLBPRIO(i));
           end generate TIEC440DCUWRURGENTPLBPRIO_DELAY;
              VitalWireDelay (TIEC440ENDIANRESET_ipd,TIEC440ENDIANRESET,tipd_TIEC440ENDIANRESET);
           TIEC440ERPNRESET_DELAY : for i in 0 to 3 generate
              VitalWireDelay (TIEC440ERPNRESET_ipd(i),TIEC440ERPNRESET(i),tipd_TIEC440ERPNRESET(i));
           end generate TIEC440ERPNRESET_DELAY;
           TIEC440ICURDFETCHPLBPRIO_DELAY : for i in 0 to 1 generate
              VitalWireDelay (TIEC440ICURDFETCHPLBPRIO_ipd(i),TIEC440ICURDFETCHPLBPRIO(i),tipd_TIEC440ICURDFETCHPLBPRIO(i));
           end generate TIEC440ICURDFETCHPLBPRIO_DELAY;
           TIEC440ICURDSPECPLBPRIO_DELAY : for i in 0 to 1 generate
              VitalWireDelay (TIEC440ICURDSPECPLBPRIO_ipd(i),TIEC440ICURDSPECPLBPRIO(i),tipd_TIEC440ICURDSPECPLBPRIO(i));
           end generate TIEC440ICURDSPECPLBPRIO_DELAY;
           TIEC440ICURDTOUCHPLBPRIO_DELAY : for i in 0 to 1 generate
              VitalWireDelay (TIEC440ICURDTOUCHPLBPRIO_ipd(i),TIEC440ICURDTOUCHPLBPRIO(i),tipd_TIEC440ICURDTOUCHPLBPRIO(i));
           end generate TIEC440ICURDTOUCHPLBPRIO_DELAY;
           TIEC440PIR_DELAY : for i in 28 to 31 generate
              VitalWireDelay (TIEC440PIR_ipd(i),TIEC440PIR(i),tipd_TIEC440PIR(i));
           end generate TIEC440PIR_DELAY;
           TIEC440PVR_DELAY : for i in 28 to 31 generate
              VitalWireDelay (TIEC440PVR_ipd(i),TIEC440PVR(i),tipd_TIEC440PVR(i));
           end generate TIEC440PVR_DELAY;
           TIEC440USERRESET_DELAY : for i in 0 to 3 generate
              VitalWireDelay (TIEC440USERRESET_ipd(i),TIEC440USERRESET(i),tipd_TIEC440USERRESET(i));
           end generate TIEC440USERRESET_DELAY;
              VitalWireDelay (TRCC440TRACEDISABLE_ipd,TRCC440TRACEDISABLE,tipd_TRCC440TRACEDISABLE);
              VitalWireDelay (TRCC440TRIGGEREVENTIN_ipd,TRCC440TRIGGEREVENTIN,tipd_TRCC440TRIGGEREVENTIN);
	end block;

	SignalDelay : block
	begin
	VitalSignalDelay (PLBPPCS0RNW_dly,PLBPPCS0RNW_ipd,tisd_PLBPPCS0RNW_CPMPPCS0PLBCLK);
	VitalSignalDelay (PLBPPCS1RNW_dly,PLBPPCS1RNW_ipd,tisd_PLBPPCS1RNW_CPMPPCS1PLBCLK);
	VitalSignalDelay (CPMINTERCONNECTCLKNTO1_dly,CPMINTERCONNECTCLKNTO1_ipd,tisd_CPMINTERCONNECTCLKNTO1_CPMINTERCONNECTCLK);
	VitalSignalDelay (DCRPPCDMACK_dly,DCRPPCDMACK_ipd,tisd_DCRPPCDMACK_CPMDCRCLK);
	DCRPPCDMDBUSIN_DELAY : for i in 0 to 31 generate
	VitalSignalDelay (DCRPPCDMDBUSIN_dly(i),DCRPPCDMDBUSIN_ipd(i),tisd_DCRPPCDMDBUSIN_CPMDCRCLK(i));
	end generate DCRPPCDMDBUSIN_DELAY;
	VitalSignalDelay (DCRPPCDMTIMEOUTWAIT_dly,DCRPPCDMTIMEOUTWAIT_ipd,tisd_DCRPPCDMTIMEOUTWAIT_CPMDCRCLK);
	VitalSignalDelay (LLDMA0RSTENGINEREQ_dly,LLDMA0RSTENGINEREQ_ipd,tisd_LLDMA0RSTENGINEREQ_CPMDMA0LLCLK);
	LLDMA0RXD_DELAY : for i in 0 to 31 generate
	VitalSignalDelay (LLDMA0RXD_dly(i),LLDMA0RXD_ipd(i),tisd_LLDMA0RXD_CPMDMA0LLCLK(i));
	end generate LLDMA0RXD_DELAY;
	VitalSignalDelay (LLDMA0RXEOFN_dly,LLDMA0RXEOFN_ipd,tisd_LLDMA0RXEOFN_CPMDMA0LLCLK);
	VitalSignalDelay (LLDMA0RXEOPN_dly,LLDMA0RXEOPN_ipd,tisd_LLDMA0RXEOPN_CPMDMA0LLCLK);
	LLDMA0RXREM_DELAY : for i in 0 to 3 generate
	VitalSignalDelay (LLDMA0RXREM_dly(i),LLDMA0RXREM_ipd(i),tisd_LLDMA0RXREM_CPMDMA0LLCLK(i));
	end generate LLDMA0RXREM_DELAY;
	VitalSignalDelay (LLDMA0RXSOFN_dly,LLDMA0RXSOFN_ipd,tisd_LLDMA0RXSOFN_CPMDMA0LLCLK);
	VitalSignalDelay (LLDMA0RXSOPN_dly,LLDMA0RXSOPN_ipd,tisd_LLDMA0RXSOPN_CPMDMA0LLCLK);
	VitalSignalDelay (LLDMA0RXSRCRDYN_dly,LLDMA0RXSRCRDYN_ipd,tisd_LLDMA0RXSRCRDYN_CPMDMA0LLCLK);
	VitalSignalDelay (LLDMA0TXDSTRDYN_dly,LLDMA0TXDSTRDYN_ipd,tisd_LLDMA0TXDSTRDYN_CPMDMA0LLCLK);
	VitalSignalDelay (LLDMA1RSTENGINEREQ_dly,LLDMA1RSTENGINEREQ_ipd,tisd_LLDMA1RSTENGINEREQ_CPMDMA1LLCLK);
	LLDMA1RXD_DELAY : for i in 0 to 31 generate
	VitalSignalDelay (LLDMA1RXD_dly(i),LLDMA1RXD_ipd(i),tisd_LLDMA1RXD_CPMDMA1LLCLK(i));
	end generate LLDMA1RXD_DELAY;
	VitalSignalDelay (LLDMA1RXEOFN_dly,LLDMA1RXEOFN_ipd,tisd_LLDMA1RXEOFN_CPMDMA1LLCLK);
	VitalSignalDelay (LLDMA1RXEOPN_dly,LLDMA1RXEOPN_ipd,tisd_LLDMA1RXEOPN_CPMDMA1LLCLK);
	LLDMA1RXREM_DELAY : for i in 0 to 3 generate
	VitalSignalDelay (LLDMA1RXREM_dly(i),LLDMA1RXREM_ipd(i),tisd_LLDMA1RXREM_CPMDMA1LLCLK(i));
	end generate LLDMA1RXREM_DELAY;
	VitalSignalDelay (LLDMA1RXSOFN_dly,LLDMA1RXSOFN_ipd,tisd_LLDMA1RXSOFN_CPMDMA1LLCLK);
	VitalSignalDelay (LLDMA1RXSOPN_dly,LLDMA1RXSOPN_ipd,tisd_LLDMA1RXSOPN_CPMDMA1LLCLK);
	VitalSignalDelay (LLDMA1RXSRCRDYN_dly,LLDMA1RXSRCRDYN_ipd,tisd_LLDMA1RXSRCRDYN_CPMDMA1LLCLK);
	VitalSignalDelay (LLDMA1TXDSTRDYN_dly,LLDMA1TXDSTRDYN_ipd,tisd_LLDMA1TXDSTRDYN_CPMDMA1LLCLK);
	VitalSignalDelay (LLDMA2RSTENGINEREQ_dly,LLDMA2RSTENGINEREQ_ipd,tisd_LLDMA2RSTENGINEREQ_CPMDMA2LLCLK);
	LLDMA2RXD_DELAY : for i in 0 to 31 generate
	VitalSignalDelay (LLDMA2RXD_dly(i),LLDMA2RXD_ipd(i),tisd_LLDMA2RXD_CPMDMA2LLCLK(i));
	end generate LLDMA2RXD_DELAY;
	VitalSignalDelay (LLDMA2RXEOFN_dly,LLDMA2RXEOFN_ipd,tisd_LLDMA2RXEOFN_CPMDMA2LLCLK);
	VitalSignalDelay (LLDMA2RXEOPN_dly,LLDMA2RXEOPN_ipd,tisd_LLDMA2RXEOPN_CPMDMA2LLCLK);
	LLDMA2RXREM_DELAY : for i in 0 to 3 generate
	VitalSignalDelay (LLDMA2RXREM_dly(i),LLDMA2RXREM_ipd(i),tisd_LLDMA2RXREM_CPMDMA2LLCLK(i));
	end generate LLDMA2RXREM_DELAY;
	VitalSignalDelay (LLDMA2RXSOFN_dly,LLDMA2RXSOFN_ipd,tisd_LLDMA2RXSOFN_CPMDMA2LLCLK);
	VitalSignalDelay (LLDMA2RXSOPN_dly,LLDMA2RXSOPN_ipd,tisd_LLDMA2RXSOPN_CPMDMA2LLCLK);
	VitalSignalDelay (LLDMA2RXSRCRDYN_dly,LLDMA2RXSRCRDYN_ipd,tisd_LLDMA2RXSRCRDYN_CPMDMA2LLCLK);
	VitalSignalDelay (LLDMA2TXDSTRDYN_dly,LLDMA2TXDSTRDYN_ipd,tisd_LLDMA2TXDSTRDYN_CPMDMA2LLCLK);
	VitalSignalDelay (LLDMA3RSTENGINEREQ_dly,LLDMA3RSTENGINEREQ_ipd,tisd_LLDMA3RSTENGINEREQ_CPMDMA3LLCLK);
	LLDMA3RXD_DELAY : for i in 0 to 31 generate
	VitalSignalDelay (LLDMA3RXD_dly(i),LLDMA3RXD_ipd(i),tisd_LLDMA3RXD_CPMDMA3LLCLK(i));
	end generate LLDMA3RXD_DELAY;
	VitalSignalDelay (LLDMA3RXEOFN_dly,LLDMA3RXEOFN_ipd,tisd_LLDMA3RXEOFN_CPMDMA3LLCLK);
	VitalSignalDelay (LLDMA3RXEOPN_dly,LLDMA3RXEOPN_ipd,tisd_LLDMA3RXEOPN_CPMDMA3LLCLK);
	LLDMA3RXREM_DELAY : for i in 0 to 3 generate
	VitalSignalDelay (LLDMA3RXREM_dly(i),LLDMA3RXREM_ipd(i),tisd_LLDMA3RXREM_CPMDMA3LLCLK(i));
	end generate LLDMA3RXREM_DELAY;
	VitalSignalDelay (LLDMA3RXSOFN_dly,LLDMA3RXSOFN_ipd,tisd_LLDMA3RXSOFN_CPMDMA3LLCLK);
	VitalSignalDelay (LLDMA3RXSOPN_dly,LLDMA3RXSOPN_ipd,tisd_LLDMA3RXSOPN_CPMDMA3LLCLK);
	VitalSignalDelay (LLDMA3RXSRCRDYN_dly,LLDMA3RXSRCRDYN_ipd,tisd_LLDMA3RXSRCRDYN_CPMDMA3LLCLK);
	VitalSignalDelay (LLDMA3TXDSTRDYN_dly,LLDMA3TXDSTRDYN_ipd,tisd_LLDMA3TXDSTRDYN_CPMDMA3LLCLK);
	VitalSignalDelay (PLBPPCMADDRACK_dly,PLBPPCMADDRACK_ipd,tisd_PLBPPCMADDRACK_CPMPPCMPLBCLK);
	VitalSignalDelay (PLBPPCMMBUSY_dly,PLBPPCMMBUSY_ipd,tisd_PLBPPCMMBUSY_CPMPPCMPLBCLK);
	VitalSignalDelay (PLBPPCMMIRQ_dly,PLBPPCMMIRQ_ipd,tisd_PLBPPCMMIRQ_CPMPPCMPLBCLK);
	VitalSignalDelay (PLBPPCMMRDERR_dly,PLBPPCMMRDERR_ipd,tisd_PLBPPCMMRDERR_CPMPPCMPLBCLK);
	VitalSignalDelay (PLBPPCMMWRERR_dly,PLBPPCMMWRERR_ipd,tisd_PLBPPCMMWRERR_CPMPPCMPLBCLK);
	VitalSignalDelay (PLBPPCMRDBTERM_dly,PLBPPCMRDBTERM_ipd,tisd_PLBPPCMRDBTERM_CPMPPCMPLBCLK);
	VitalSignalDelay (PLBPPCMRDDACK_dly,PLBPPCMRDDACK_ipd,tisd_PLBPPCMRDDACK_CPMPPCMPLBCLK);
	PLBPPCMRDDBUS_DELAY : for i in 0 to 127 generate
	VitalSignalDelay (PLBPPCMRDDBUS_dly(i),PLBPPCMRDDBUS_ipd(i),tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(i));
	end generate PLBPPCMRDDBUS_DELAY;
	PLBPPCMRDPENDPRI_DELAY : for i in 0 to 1 generate
	VitalSignalDelay (PLBPPCMRDPENDPRI_dly(i),PLBPPCMRDPENDPRI_ipd(i),tisd_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK(i));
	end generate PLBPPCMRDPENDPRI_DELAY;
	VitalSignalDelay (PLBPPCMRDPENDREQ_dly,PLBPPCMRDPENDREQ_ipd,tisd_PLBPPCMRDPENDREQ_CPMPPCMPLBCLK);
	PLBPPCMRDWDADDR_DELAY : for i in 0 to 3 generate
	VitalSignalDelay (PLBPPCMRDWDADDR_dly(i),PLBPPCMRDWDADDR_ipd(i),tisd_PLBPPCMRDWDADDR_CPMPPCMPLBCLK(i));
	end generate PLBPPCMRDWDADDR_DELAY;
	VitalSignalDelay (PLBPPCMREARBITRATE_dly,PLBPPCMREARBITRATE_ipd,tisd_PLBPPCMREARBITRATE_CPMPPCMPLBCLK);
	PLBPPCMREQPRI_DELAY : for i in 0 to 1 generate
	VitalSignalDelay (PLBPPCMREQPRI_dly(i),PLBPPCMREQPRI_ipd(i),tisd_PLBPPCMREQPRI_CPMPPCMPLBCLK(i));
	end generate PLBPPCMREQPRI_DELAY;
	PLBPPCMSSIZE_DELAY : for i in 0 to 1 generate
	VitalSignalDelay (PLBPPCMSSIZE_dly(i),PLBPPCMSSIZE_ipd(i),tisd_PLBPPCMSSIZE_CPMPPCMPLBCLK(i));
	end generate PLBPPCMSSIZE_DELAY;
	VitalSignalDelay (PLBPPCMTIMEOUT_dly,PLBPPCMTIMEOUT_ipd,tisd_PLBPPCMTIMEOUT_CPMPPCMPLBCLK);
	VitalSignalDelay (PLBPPCMWRBTERM_dly,PLBPPCMWRBTERM_ipd,tisd_PLBPPCMWRBTERM_CPMPPCMPLBCLK);
	VitalSignalDelay (PLBPPCMWRDACK_dly,PLBPPCMWRDACK_ipd,tisd_PLBPPCMWRDACK_CPMPPCMPLBCLK);
	PLBPPCMWRPENDPRI_DELAY : for i in 0 to 1 generate
	VitalSignalDelay (PLBPPCMWRPENDPRI_dly(i),PLBPPCMWRPENDPRI_ipd(i),tisd_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK(i));
	end generate PLBPPCMWRPENDPRI_DELAY;
	VitalSignalDelay (PLBPPCMWRPENDREQ_dly,PLBPPCMWRPENDREQ_ipd,tisd_PLBPPCMWRPENDREQ_CPMPPCMPLBCLK);
	VitalSignalDelay (PLBPPCS0ABORT_dly,PLBPPCS0ABORT_ipd,tisd_PLBPPCS0ABORT_CPMPPCS0PLBCLK);
	PLBPPCS0ABUS_DELAY : for i in 0 to 31 generate
	VitalSignalDelay (PLBPPCS0ABUS_dly(i),PLBPPCS0ABUS_ipd(i),tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(i));
	end generate PLBPPCS0ABUS_DELAY;
	PLBPPCS0BE_DELAY : for i in 0 to 15 generate
	VitalSignalDelay (PLBPPCS0BE_dly(i),PLBPPCS0BE_ipd(i),tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(i));
	end generate PLBPPCS0BE_DELAY;
	VitalSignalDelay (PLBPPCS0BUSLOCK_dly,PLBPPCS0BUSLOCK_ipd,tisd_PLBPPCS0BUSLOCK_CPMPPCS0PLBCLK);
	VitalSignalDelay (PLBPPCS0LOCKERR_dly,PLBPPCS0LOCKERR_ipd,tisd_PLBPPCS0LOCKERR_CPMPPCS0PLBCLK);
	PLBPPCS0MASTERID_DELAY : for i in 0 to 1 generate
	VitalSignalDelay (PLBPPCS0MASTERID_dly(i),PLBPPCS0MASTERID_ipd(i),tisd_PLBPPCS0MASTERID_CPMPPCS0PLBCLK(i));
	end generate PLBPPCS0MASTERID_DELAY;
	PLBPPCS0MSIZE_DELAY : for i in 0 to 1 generate
	VitalSignalDelay (PLBPPCS0MSIZE_dly(i),PLBPPCS0MSIZE_ipd(i),tisd_PLBPPCS0MSIZE_CPMPPCS0PLBCLK(i));
	end generate PLBPPCS0MSIZE_DELAY;
	VitalSignalDelay (PLBPPCS0PAVALID_dly,PLBPPCS0PAVALID_ipd,tisd_PLBPPCS0PAVALID_CPMPPCS0PLBCLK);
	VitalSignalDelay (PLBPPCS0RDBURST_dly,PLBPPCS0RDBURST_ipd,tisd_PLBPPCS0RDBURST_CPMPPCS0PLBCLK);
	PLBPPCS0RDPENDPRI_DELAY : for i in 0 to 1 generate
	VitalSignalDelay (PLBPPCS0RDPENDPRI_dly(i),PLBPPCS0RDPENDPRI_ipd(i),tisd_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK(i));
	end generate PLBPPCS0RDPENDPRI_DELAY;
	VitalSignalDelay (PLBPPCS0RDPENDREQ_dly,PLBPPCS0RDPENDREQ_ipd,tisd_PLBPPCS0RDPENDREQ_CPMPPCS0PLBCLK);
	VitalSignalDelay (PLBPPCS0RDPRIM_dly,PLBPPCS0RDPRIM_ipd,tisd_PLBPPCS0RDPRIM_CPMPPCS0PLBCLK);
	PLBPPCS0REQPRI_DELAY : for i in 0 to 1 generate
	VitalSignalDelay (PLBPPCS0REQPRI_dly(i),PLBPPCS0REQPRI_ipd(i),tisd_PLBPPCS0REQPRI_CPMPPCS0PLBCLK(i));
	end generate PLBPPCS0REQPRI_DELAY;
	VitalSignalDelay (PLBPPCS0SAVALID_dly,PLBPPCS0SAVALID_ipd,tisd_PLBPPCS0SAVALID_CPMPPCS0PLBCLK);
	PLBPPCS0SIZE_DELAY : for i in 0 to 3 generate
	VitalSignalDelay (PLBPPCS0SIZE_dly(i),PLBPPCS0SIZE_ipd(i),tisd_PLBPPCS0SIZE_CPMPPCS0PLBCLK(i));
	end generate PLBPPCS0SIZE_DELAY;
	PLBPPCS0TATTRIBUTE_DELAY : for i in 0 to 15 generate
	VitalSignalDelay (PLBPPCS0TATTRIBUTE_dly(i),PLBPPCS0TATTRIBUTE_ipd(i),tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(i));
	end generate PLBPPCS0TATTRIBUTE_DELAY;
	PLBPPCS0TYPE_DELAY : for i in 0 to 2 generate
	VitalSignalDelay (PLBPPCS0TYPE_dly(i),PLBPPCS0TYPE_ipd(i),tisd_PLBPPCS0TYPE_CPMPPCS0PLBCLK(i));
	end generate PLBPPCS0TYPE_DELAY;
	PLBPPCS0UABUS_DELAY : for i in 28 to 31 generate
	VitalSignalDelay (PLBPPCS0UABUS_dly(i),PLBPPCS0UABUS_ipd(i),tisd_PLBPPCS0UABUS_CPMPPCS0PLBCLK(i));
	end generate PLBPPCS0UABUS_DELAY;
	VitalSignalDelay (PLBPPCS0WRBURST_dly,PLBPPCS0WRBURST_ipd,tisd_PLBPPCS0WRBURST_CPMPPCS0PLBCLK);
	PLBPPCS0WRDBUS_DELAY : for i in 0 to 127 generate
	VitalSignalDelay (PLBPPCS0WRDBUS_dly(i),PLBPPCS0WRDBUS_ipd(i),tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(i));
	end generate PLBPPCS0WRDBUS_DELAY;
	PLBPPCS0WRPENDPRI_DELAY : for i in 0 to 1 generate
	VitalSignalDelay (PLBPPCS0WRPENDPRI_dly(i),PLBPPCS0WRPENDPRI_ipd(i),tisd_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK(i));
	end generate PLBPPCS0WRPENDPRI_DELAY;
	VitalSignalDelay (PLBPPCS0WRPENDREQ_dly,PLBPPCS0WRPENDREQ_ipd,tisd_PLBPPCS0WRPENDREQ_CPMPPCS0PLBCLK);
	VitalSignalDelay (PLBPPCS0WRPRIM_dly,PLBPPCS0WRPRIM_ipd,tisd_PLBPPCS0WRPRIM_CPMPPCS0PLBCLK);
	VitalSignalDelay (PLBPPCS1ABORT_dly,PLBPPCS1ABORT_ipd,tisd_PLBPPCS1ABORT_CPMPPCS1PLBCLK);
	PLBPPCS1ABUS_DELAY : for i in 0 to 31 generate
	VitalSignalDelay (PLBPPCS1ABUS_dly(i),PLBPPCS1ABUS_ipd(i),tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(i));
	end generate PLBPPCS1ABUS_DELAY;
	PLBPPCS1BE_DELAY : for i in 0 to 15 generate
	VitalSignalDelay (PLBPPCS1BE_dly(i),PLBPPCS1BE_ipd(i),tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(i));
	end generate PLBPPCS1BE_DELAY;
	VitalSignalDelay (PLBPPCS1BUSLOCK_dly,PLBPPCS1BUSLOCK_ipd,tisd_PLBPPCS1BUSLOCK_CPMPPCS1PLBCLK);
	VitalSignalDelay (PLBPPCS1LOCKERR_dly,PLBPPCS1LOCKERR_ipd,tisd_PLBPPCS1LOCKERR_CPMPPCS1PLBCLK);
	PLBPPCS1MASTERID_DELAY : for i in 0 to 1 generate
	VitalSignalDelay (PLBPPCS1MASTERID_dly(i),PLBPPCS1MASTERID_ipd(i),tisd_PLBPPCS1MASTERID_CPMPPCS1PLBCLK(i));
	end generate PLBPPCS1MASTERID_DELAY;
	PLBPPCS1MSIZE_DELAY : for i in 0 to 1 generate
	VitalSignalDelay (PLBPPCS1MSIZE_dly(i),PLBPPCS1MSIZE_ipd(i),tisd_PLBPPCS1MSIZE_CPMPPCS1PLBCLK(i));
	end generate PLBPPCS1MSIZE_DELAY;
	VitalSignalDelay (PLBPPCS1PAVALID_dly,PLBPPCS1PAVALID_ipd,tisd_PLBPPCS1PAVALID_CPMPPCS1PLBCLK);
	VitalSignalDelay (PLBPPCS1RDBURST_dly,PLBPPCS1RDBURST_ipd,tisd_PLBPPCS1RDBURST_CPMPPCS1PLBCLK);
	PLBPPCS1RDPENDPRI_DELAY : for i in 0 to 1 generate
	VitalSignalDelay (PLBPPCS1RDPENDPRI_dly(i),PLBPPCS1RDPENDPRI_ipd(i),tisd_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK(i));
	end generate PLBPPCS1RDPENDPRI_DELAY;
	VitalSignalDelay (PLBPPCS1RDPENDREQ_dly,PLBPPCS1RDPENDREQ_ipd,tisd_PLBPPCS1RDPENDREQ_CPMPPCS1PLBCLK);
	VitalSignalDelay (PLBPPCS1RDPRIM_dly,PLBPPCS1RDPRIM_ipd,tisd_PLBPPCS1RDPRIM_CPMPPCS1PLBCLK);
	PLBPPCS1REQPRI_DELAY : for i in 0 to 1 generate
	VitalSignalDelay (PLBPPCS1REQPRI_dly(i),PLBPPCS1REQPRI_ipd(i),tisd_PLBPPCS1REQPRI_CPMPPCS1PLBCLK(i));
	end generate PLBPPCS1REQPRI_DELAY;
	VitalSignalDelay (PLBPPCS1SAVALID_dly,PLBPPCS1SAVALID_ipd,tisd_PLBPPCS1SAVALID_CPMPPCS1PLBCLK);
	PLBPPCS1SIZE_DELAY : for i in 0 to 3 generate
	VitalSignalDelay (PLBPPCS1SIZE_dly(i),PLBPPCS1SIZE_ipd(i),tisd_PLBPPCS1SIZE_CPMPPCS1PLBCLK(i));
	end generate PLBPPCS1SIZE_DELAY;
	PLBPPCS1TATTRIBUTE_DELAY : for i in 0 to 15 generate
	VitalSignalDelay (PLBPPCS1TATTRIBUTE_dly(i),PLBPPCS1TATTRIBUTE_ipd(i),tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(i));
	end generate PLBPPCS1TATTRIBUTE_DELAY;
	PLBPPCS1TYPE_DELAY : for i in 0 to 2 generate
	VitalSignalDelay (PLBPPCS1TYPE_dly(i),PLBPPCS1TYPE_ipd(i),tisd_PLBPPCS1TYPE_CPMPPCS1PLBCLK(i));
	end generate PLBPPCS1TYPE_DELAY;
	PLBPPCS1UABUS_DELAY : for i in 28 to 31 generate
	VitalSignalDelay (PLBPPCS1UABUS_dly(i),PLBPPCS1UABUS_ipd(i),tisd_PLBPPCS1UABUS_CPMPPCS1PLBCLK(i));
	end generate PLBPPCS1UABUS_DELAY;
	VitalSignalDelay (PLBPPCS1WRBURST_dly,PLBPPCS1WRBURST_ipd,tisd_PLBPPCS1WRBURST_CPMPPCS1PLBCLK);
	PLBPPCS1WRDBUS_DELAY : for i in 0 to 127 generate
	VitalSignalDelay (PLBPPCS1WRDBUS_dly(i),PLBPPCS1WRDBUS_ipd(i),tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(i));
	end generate PLBPPCS1WRDBUS_DELAY;
	PLBPPCS1WRPENDPRI_DELAY : for i in 0 to 1 generate
	VitalSignalDelay (PLBPPCS1WRPENDPRI_dly(i),PLBPPCS1WRPENDPRI_ipd(i),tisd_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK(i));
	end generate PLBPPCS1WRPENDPRI_DELAY;
	VitalSignalDelay (PLBPPCS1WRPENDREQ_dly,PLBPPCS1WRPENDREQ_ipd,tisd_PLBPPCS1WRPENDREQ_CPMPPCS1PLBCLK);
	VitalSignalDelay (PLBPPCS1WRPRIM_dly,PLBPPCS1WRPRIM_ipd,tisd_PLBPPCS1WRPRIM_CPMPPCS1PLBCLK);
	VitalSignalDelay (CPMC440CORECLOCKINACTIVE_dly,CPMC440CORECLOCKINACTIVE_ipd,tisd_CPMC440CORECLOCKINACTIVE_JTGC440TCK);
	VitalSignalDelay (DBGC440DEBUGHALT_dly,DBGC440DEBUGHALT_ipd,tisd_DBGC440DEBUGHALT_CPMC440CLK);
	DBGC440SYSTEMSTATUS_DELAY : for i in 0 to 4 generate
	VitalSignalDelay (DBGC440SYSTEMSTATUS_dly(i),DBGC440SYSTEMSTATUS_ipd(i),tisd_DBGC440SYSTEMSTATUS_JTGC440TCK(i));
	end generate DBGC440SYSTEMSTATUS_DELAY;
	VitalSignalDelay (DBGC440UNCONDDEBUGEVENT_dly,DBGC440UNCONDDEBUGEVENT_ipd,tisd_DBGC440UNCONDDEBUGEVENT_CPMC440CLK);
	DCRPPCDSABUS_DELAY : for i in 0 to 9 generate
	VitalSignalDelay (DCRPPCDSABUS_dly(i),DCRPPCDSABUS_ipd(i),tisd_DCRPPCDSABUS_CPMDCRCLK(i));
	end generate DCRPPCDSABUS_DELAY;
	DCRPPCDSDBUSOUT_DELAY : for i in 0 to 31 generate
	VitalSignalDelay (DCRPPCDSDBUSOUT_dly(i),DCRPPCDSDBUSOUT_ipd(i),tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(i));
	end generate DCRPPCDSDBUSOUT_DELAY;
	VitalSignalDelay (DCRPPCDSREAD_dly,DCRPPCDSREAD_ipd,tisd_DCRPPCDSREAD_CPMDCRCLK);
	VitalSignalDelay (DCRPPCDSWRITE_dly,DCRPPCDSWRITE_ipd,tisd_DCRPPCDSWRITE_CPMDCRCLK);
	VitalSignalDelay (FCMAPUCONFIRMINSTR_dly,FCMAPUCONFIRMINSTR_ipd,tisd_FCMAPUCONFIRMINSTR_CPMFCMCLK);
	FCMAPUCR_DELAY : for i in 0 to 3 generate
	VitalSignalDelay (FCMAPUCR_dly(i),FCMAPUCR_ipd(i),tisd_FCMAPUCR_CPMFCMCLK(i));
	end generate FCMAPUCR_DELAY;
	VitalSignalDelay (FCMAPUDONE_dly,FCMAPUDONE_ipd,tisd_FCMAPUDONE_CPMFCMCLK);
	VitalSignalDelay (FCMAPUEXCEPTION_dly,FCMAPUEXCEPTION_ipd,tisd_FCMAPUEXCEPTION_CPMFCMCLK);
	VitalSignalDelay (FCMAPUFPSCRFEX_dly,FCMAPUFPSCRFEX_ipd,tisd_FCMAPUFPSCRFEX_CPMFCMCLK);
	FCMAPURESULT_DELAY : for i in 0 to 31 generate
	VitalSignalDelay (FCMAPURESULT_dly(i),FCMAPURESULT_ipd(i),tisd_FCMAPURESULT_CPMFCMCLK(i));
	end generate FCMAPURESULT_DELAY;
	VitalSignalDelay (FCMAPURESULTVALID_dly,FCMAPURESULTVALID_ipd,tisd_FCMAPURESULTVALID_CPMFCMCLK);
	VitalSignalDelay (FCMAPUSLEEPNOTREADY_dly,FCMAPUSLEEPNOTREADY_ipd,tisd_FCMAPUSLEEPNOTREADY_CPMFCMCLK);
	FCMAPUSTOREDATA_DELAY : for i in 0 to 127 generate
	VitalSignalDelay (FCMAPUSTOREDATA_dly(i),FCMAPUSTOREDATA_ipd(i),tisd_FCMAPUSTOREDATA_CPMFCMCLK(i));
	end generate FCMAPUSTOREDATA_DELAY;
	VitalSignalDelay (JTGC440TDI_dly,JTGC440TDI_ipd,tisd_JTGC440TDI_JTGC440TCK);
	VitalSignalDelay (JTGC440TMS_dly,JTGC440TMS_ipd,tisd_JTGC440TMS_JTGC440TCK);
	VitalSignalDelay (MCMIADDRREADYTOACCEPT_dly,MCMIADDRREADYTOACCEPT_ipd,tisd_MCMIADDRREADYTOACCEPT_CPMMCCLK);
	MCMIREADDATA_DELAY : for i in 0 to 127 generate
	VitalSignalDelay (MCMIREADDATA_dly(i),MCMIREADDATA_ipd(i),tisd_MCMIREADDATA_CPMMCCLK(i));
	end generate MCMIREADDATA_DELAY;
	VitalSignalDelay (MCMIREADDATAERR_dly,MCMIREADDATAERR_ipd,tisd_MCMIREADDATAERR_CPMMCCLK);
	VitalSignalDelay (MCMIREADDATAVALID_dly,MCMIREADDATAVALID_ipd,tisd_MCMIREADDATAVALID_CPMMCCLK);
	VitalSignalDelay (TRCC440TRACEDISABLE_dly,TRCC440TRACEDISABLE_ipd,tisd_TRCC440TRACEDISABLE_CPMC440CLK);
	VitalSignalDelay (TRCC440TRIGGEREVENTIN_dly,TRCC440TRIGGEREVENTIN_ipd,tisd_TRCC440TRIGGEREVENTIN_CPMC440CLK);

	VitalSignalDelay (CPMPPCS0PLBCLK_dly,CPMPPCS0PLBCLK_ipd,ticd_CPMPPCS0PLBCLK);
	VitalSignalDelay (CPMPPCS1PLBCLK_dly,CPMPPCS1PLBCLK_ipd,ticd_CPMPPCS1PLBCLK);
	VitalSignalDelay (CPMINTERCONNECTCLK_dly,CPMINTERCONNECTCLK_ipd,ticd_CPMINTERCONNECTCLK);
	VitalSignalDelay (CPMDCRCLK_dly,CPMDCRCLK_ipd,ticd_CPMDCRCLK);
	VitalSignalDelay (CPMDMA0LLCLK_dly,CPMDMA0LLCLK_ipd,ticd_CPMDMA0LLCLK);
	VitalSignalDelay (CPMDMA1LLCLK_dly,CPMDMA1LLCLK_ipd,ticd_CPMDMA1LLCLK);
	VitalSignalDelay (CPMDMA2LLCLK_dly,CPMDMA2LLCLK_ipd,ticd_CPMDMA2LLCLK);
	VitalSignalDelay (CPMDMA3LLCLK_dly,CPMDMA3LLCLK_ipd,ticd_CPMDMA3LLCLK);
	VitalSignalDelay (CPMPPCMPLBCLK_dly,CPMPPCMPLBCLK_ipd,ticd_CPMPPCMPLBCLK);
	VitalSignalDelay (JTGC440TCK_dly,JTGC440TCK_ipd,ticd_JTGC440TCK);
	VitalSignalDelay (CPMC440CLK_dly,CPMC440CLK_ipd,ticd_CPMC440CLK);
	VitalSignalDelay (CPMFCMCLK_dly,CPMFCMCLK_ipd,ticd_CPMFCMCLK);
	VitalSignalDelay (CPMMCCLK_dly,CPMMCCLK_ipd,ticd_CPMMCCLK);
	end block;

	CPMC440CLKEN_dly <= CPMC440CLKEN_ipd;
	CPMINTERCONNECTCLKEN_dly <= CPMINTERCONNECTCLKEN_ipd;
	EICC440CRITIRQ_dly <= EICC440CRITIRQ_ipd;
	EICC440EXTIRQ_dly <= EICC440EXTIRQ_ipd;
	JTGC440TRSTNEG_dly <= JTGC440TRSTNEG_ipd;
	RSTC440RESETCHIP_dly <= RSTC440RESETCHIP_ipd;
	RSTC440RESETCORE_dly <= RSTC440RESETCORE_ipd;
	RSTC440RESETSYSTEM_dly <= RSTC440RESETSYSTEM_ipd;
	TIEC440DCURDLDCACHEPLBPRIO_dly <= TIEC440DCURDLDCACHEPLBPRIO_ipd;
	TIEC440DCURDNONCACHEPLBPRIO_dly <= TIEC440DCURDNONCACHEPLBPRIO_ipd;
	TIEC440DCURDTOUCHPLBPRIO_dly <= TIEC440DCURDTOUCHPLBPRIO_ipd;
	TIEC440DCURDURGENTPLBPRIO_dly <= TIEC440DCURDURGENTPLBPRIO_ipd;
	TIEC440DCUWRFLUSHPLBPRIO_dly <= TIEC440DCUWRFLUSHPLBPRIO_ipd;
	TIEC440DCUWRSTOREPLBPRIO_dly <= TIEC440DCUWRSTOREPLBPRIO_ipd;
	TIEC440DCUWRURGENTPLBPRIO_dly <= TIEC440DCUWRURGENTPLBPRIO_ipd;
	TIEC440ENDIANRESET_dly <= TIEC440ENDIANRESET_ipd;
	TIEC440ERPNRESET_dly <= TIEC440ERPNRESET_ipd;
	TIEC440ICURDFETCHPLBPRIO_dly <= TIEC440ICURDFETCHPLBPRIO_ipd;
	TIEC440ICURDSPECPLBPRIO_dly <= TIEC440ICURDSPECPLBPRIO_ipd;
	TIEC440ICURDTOUCHPLBPRIO_dly <= TIEC440ICURDTOUCHPLBPRIO_ipd;
	TIEC440PIR_dly <= TIEC440PIR_ipd;
	TIEC440PVR_dly <= TIEC440PVR_ipd;
	TIEC440USERRESET_dly <= TIEC440USERRESET_ipd;
	TIEDCRBASEADDR_dly <= TIEDCRBASEADDR_ipd;

	APUFCMDECFPUOP_out <= APUFCMDECFPUOP_outdelay after OUT_DELAY;
	APUFCMDECLDSTXFERSIZE_out <= APUFCMDECLDSTXFERSIZE_outdelay after OUT_DELAY;
	APUFCMDECLOAD_out <= APUFCMDECLOAD_outdelay after OUT_DELAY;
	APUFCMDECNONAUTON_out <= APUFCMDECNONAUTON_outdelay after OUT_DELAY;
	APUFCMDECSTORE_out <= APUFCMDECSTORE_outdelay after OUT_DELAY;
	APUFCMDECUDIVALID_out <= APUFCMDECUDIVALID_outdelay after OUT_DELAY;
	APUFCMDECUDI_out <= APUFCMDECUDI_outdelay after OUT_DELAY;
	APUFCMENDIAN_out <= APUFCMENDIAN_outdelay after OUT_DELAY;
	APUFCMFLUSH_out <= APUFCMFLUSH_outdelay after OUT_DELAY;
	APUFCMINSTRUCTION_out <= APUFCMINSTRUCTION_outdelay after OUT_DELAY;
	APUFCMINSTRVALID_out <= APUFCMINSTRVALID_outdelay after OUT_DELAY;
	APUFCMLOADBYTEADDR_out <= APUFCMLOADBYTEADDR_outdelay after OUT_DELAY;
	APUFCMLOADDATA_out <= APUFCMLOADDATA_outdelay after OUT_DELAY;
	APUFCMLOADDVALID_out <= APUFCMLOADDVALID_outdelay after OUT_DELAY;
	APUFCMMSRFE0_out <= APUFCMMSRFE0_outdelay after OUT_DELAY;
	APUFCMMSRFE1_out <= APUFCMMSRFE1_outdelay after OUT_DELAY;
	APUFCMNEXTINSTRREADY_out <= APUFCMNEXTINSTRREADY_outdelay after OUT_DELAY;
	APUFCMOPERANDVALID_out <= APUFCMOPERANDVALID_outdelay after OUT_DELAY;
	APUFCMRADATA_out <= APUFCMRADATA_outdelay after OUT_DELAY;
	APUFCMRBDATA_out <= APUFCMRBDATA_outdelay after OUT_DELAY;
	APUFCMWRITEBACKOK_out <= APUFCMWRITEBACKOK_outdelay after OUT_DELAY;
	C440CPMCORESLEEPREQ_out <= C440CPMCORESLEEPREQ_outdelay after OUT_DELAY;
	C440CPMDECIRPTREQ_out <= C440CPMDECIRPTREQ_outdelay after OUT_DELAY;
	C440CPMFITIRPTREQ_out <= C440CPMFITIRPTREQ_outdelay after OUT_DELAY;
	C440CPMMSRCE_out <= C440CPMMSRCE_outdelay after OUT_DELAY;
	C440CPMMSREE_out <= C440CPMMSREE_outdelay after OUT_DELAY;
	C440CPMTIMERRESETREQ_out <= C440CPMTIMERRESETREQ_outdelay after OUT_DELAY;
	C440CPMWDIRPTREQ_out <= C440CPMWDIRPTREQ_outdelay after OUT_DELAY;
	C440DBGSYSTEMCONTROL_out <= C440DBGSYSTEMCONTROL_outdelay after OUT_DELAY;
	C440JTGTDOEN_out <= C440JTGTDOEN_outdelay after OUT_DELAY;
	C440JTGTDO_out <= C440JTGTDO_outdelay after OUT_DELAY;
	C440MACHINECHECK_out <= C440MACHINECHECK_outdelay after OUT_DELAY;
	C440RSTCHIPRESETREQ_out <= C440RSTCHIPRESETREQ_outdelay after OUT_DELAY;
	C440RSTCORERESETREQ_out <= C440RSTCORERESETREQ_outdelay after OUT_DELAY;
	C440RSTSYSTEMRESETREQ_out <= C440RSTSYSTEMRESETREQ_outdelay after OUT_DELAY;
	C440TRCBRANCHSTATUS_out <= C440TRCBRANCHSTATUS_outdelay after OUT_DELAY;
	C440TRCCYCLE_out <= C440TRCCYCLE_outdelay after OUT_DELAY;
	C440TRCEXECUTIONSTATUS_out <= C440TRCEXECUTIONSTATUS_outdelay after OUT_DELAY;
	C440TRCTRACESTATUS_out <= C440TRCTRACESTATUS_outdelay after OUT_DELAY;
	C440TRCTRIGGEREVENTOUT_out <= C440TRCTRIGGEREVENTOUT_outdelay after OUT_DELAY;
	C440TRCTRIGGEREVENTTYPE_out <= C440TRCTRIGGEREVENTTYPE_outdelay after OUT_DELAY;
	DMA0LLRSTENGINEACK_out <= DMA0LLRSTENGINEACK_outdelay after OUT_DELAY;
	DMA0LLRXDSTRDYN_out <= DMA0LLRXDSTRDYN_outdelay after OUT_DELAY;
	DMA0LLTXD_out <= DMA0LLTXD_outdelay after OUT_DELAY;
	DMA0LLTXEOFN_out <= DMA0LLTXEOFN_outdelay after OUT_DELAY;
	DMA0LLTXEOPN_out <= DMA0LLTXEOPN_outdelay after OUT_DELAY;
	DMA0LLTXREM_out <= DMA0LLTXREM_outdelay after OUT_DELAY;
	DMA0LLTXSOFN_out <= DMA0LLTXSOFN_outdelay after OUT_DELAY;
	DMA0LLTXSOPN_out <= DMA0LLTXSOPN_outdelay after OUT_DELAY;
	DMA0LLTXSRCRDYN_out <= DMA0LLTXSRCRDYN_outdelay after OUT_DELAY;
	DMA0RXIRQ_out <= DMA0RXIRQ_outdelay after OUT_DELAY;
	DMA0TXIRQ_out <= DMA0TXIRQ_outdelay after OUT_DELAY;
	DMA1LLRSTENGINEACK_out <= DMA1LLRSTENGINEACK_outdelay after OUT_DELAY;
	DMA1LLRXDSTRDYN_out <= DMA1LLRXDSTRDYN_outdelay after OUT_DELAY;
	DMA1LLTXD_out <= DMA1LLTXD_outdelay after OUT_DELAY;
	DMA1LLTXEOFN_out <= DMA1LLTXEOFN_outdelay after OUT_DELAY;
	DMA1LLTXEOPN_out <= DMA1LLTXEOPN_outdelay after OUT_DELAY;
	DMA1LLTXREM_out <= DMA1LLTXREM_outdelay after OUT_DELAY;
	DMA1LLTXSOFN_out <= DMA1LLTXSOFN_outdelay after OUT_DELAY;
	DMA1LLTXSOPN_out <= DMA1LLTXSOPN_outdelay after OUT_DELAY;
	DMA1LLTXSRCRDYN_out <= DMA1LLTXSRCRDYN_outdelay after OUT_DELAY;
	DMA1RXIRQ_out <= DMA1RXIRQ_outdelay after OUT_DELAY;
	DMA1TXIRQ_out <= DMA1TXIRQ_outdelay after OUT_DELAY;
	DMA2LLRSTENGINEACK_out <= DMA2LLRSTENGINEACK_outdelay after OUT_DELAY;
	DMA2LLRXDSTRDYN_out <= DMA2LLRXDSTRDYN_outdelay after OUT_DELAY;
	DMA2LLTXD_out <= DMA2LLTXD_outdelay after OUT_DELAY;
	DMA2LLTXEOFN_out <= DMA2LLTXEOFN_outdelay after OUT_DELAY;
	DMA2LLTXEOPN_out <= DMA2LLTXEOPN_outdelay after OUT_DELAY;
	DMA2LLTXREM_out <= DMA2LLTXREM_outdelay after OUT_DELAY;
	DMA2LLTXSOFN_out <= DMA2LLTXSOFN_outdelay after OUT_DELAY;
	DMA2LLTXSOPN_out <= DMA2LLTXSOPN_outdelay after OUT_DELAY;
	DMA2LLTXSRCRDYN_out <= DMA2LLTXSRCRDYN_outdelay after OUT_DELAY;
	DMA2RXIRQ_out <= DMA2RXIRQ_outdelay after OUT_DELAY;
	DMA2TXIRQ_out <= DMA2TXIRQ_outdelay after OUT_DELAY;
	DMA3LLRSTENGINEACK_out <= DMA3LLRSTENGINEACK_outdelay after OUT_DELAY;
	DMA3LLRXDSTRDYN_out <= DMA3LLRXDSTRDYN_outdelay after OUT_DELAY;
	DMA3LLTXD_out <= DMA3LLTXD_outdelay after OUT_DELAY;
	DMA3LLTXEOFN_out <= DMA3LLTXEOFN_outdelay after OUT_DELAY;
	DMA3LLTXEOPN_out <= DMA3LLTXEOPN_outdelay after OUT_DELAY;
	DMA3LLTXREM_out <= DMA3LLTXREM_outdelay after OUT_DELAY;
	DMA3LLTXSOFN_out <= DMA3LLTXSOFN_outdelay after OUT_DELAY;
	DMA3LLTXSOPN_out <= DMA3LLTXSOPN_outdelay after OUT_DELAY;
	DMA3LLTXSRCRDYN_out <= DMA3LLTXSRCRDYN_outdelay after OUT_DELAY;
	DMA3RXIRQ_out <= DMA3RXIRQ_outdelay after OUT_DELAY;
	DMA3TXIRQ_out <= DMA3TXIRQ_outdelay after OUT_DELAY;
	MIMCADDRESSVALID_out <= MIMCADDRESSVALID_outdelay after OUT_DELAY;
	MIMCADDRESS_out <= MIMCADDRESS_outdelay after OUT_DELAY;
	MIMCBANKCONFLICT_out <= MIMCBANKCONFLICT_outdelay after OUT_DELAY;
	MIMCBYTEENABLE_out <= MIMCBYTEENABLE_outdelay after OUT_DELAY;
	MIMCREADNOTWRITE_out <= MIMCREADNOTWRITE_outdelay after OUT_DELAY;
	MIMCROWCONFLICT_out <= MIMCROWCONFLICT_outdelay after OUT_DELAY;
	MIMCWRITEDATAVALID_out <= MIMCWRITEDATAVALID_outdelay after OUT_DELAY;
	MIMCWRITEDATA_out <= MIMCWRITEDATA_outdelay after OUT_DELAY;
	PPCCPMINTERCONNECTBUSY_out <= PPCCPMINTERCONNECTBUSY_outdelay after OUT_DELAY;
	PPCDMDCRABUS_out <= PPCDMDCRABUS_outdelay after OUT_DELAY;
	PPCDMDCRDBUSOUT_out <= PPCDMDCRDBUSOUT_outdelay after OUT_DELAY;
	PPCDMDCRREAD_out <= PPCDMDCRREAD_outdelay after OUT_DELAY;
	PPCDMDCRUABUS_out <= PPCDMDCRUABUS_outdelay after OUT_DELAY;
	PPCDMDCRWRITE_out <= PPCDMDCRWRITE_outdelay after OUT_DELAY;
	PPCDSDCRACK_out <= PPCDSDCRACK_outdelay after OUT_DELAY;
	PPCDSDCRDBUSIN_out <= PPCDSDCRDBUSIN_outdelay after OUT_DELAY;
	PPCDSDCRTIMEOUTWAIT_out <= PPCDSDCRTIMEOUTWAIT_outdelay after OUT_DELAY;
	PPCEICINTERCONNECTIRQ_out <= PPCEICINTERCONNECTIRQ_outdelay after OUT_DELAY;
	PPCMPLBABORT_out <= PPCMPLBABORT_outdelay after OUT_DELAY;
	PPCMPLBABUS_out <= PPCMPLBABUS_outdelay after OUT_DELAY;
	PPCMPLBBE_out <= PPCMPLBBE_outdelay after OUT_DELAY;
	PPCMPLBBUSLOCK_out <= PPCMPLBBUSLOCK_outdelay after OUT_DELAY;
	PPCMPLBLOCKERR_out <= PPCMPLBLOCKERR_outdelay after OUT_DELAY;
	PPCMPLBPRIORITY_out <= PPCMPLBPRIORITY_outdelay after OUT_DELAY;
	PPCMPLBRDBURST_out <= PPCMPLBRDBURST_outdelay after OUT_DELAY;
	PPCMPLBREQUEST_out <= PPCMPLBREQUEST_outdelay after OUT_DELAY;
	PPCMPLBRNW_out <= PPCMPLBRNW_outdelay after OUT_DELAY;
	PPCMPLBSIZE_out <= PPCMPLBSIZE_outdelay after OUT_DELAY;
	PPCMPLBTATTRIBUTE_out <= PPCMPLBTATTRIBUTE_outdelay after OUT_DELAY;
	PPCMPLBTYPE_out <= PPCMPLBTYPE_outdelay after OUT_DELAY;
	PPCMPLBUABUS_out <= PPCMPLBUABUS_outdelay after OUT_DELAY;
	PPCMPLBWRBURST_out <= PPCMPLBWRBURST_outdelay after OUT_DELAY;
	PPCMPLBWRDBUS_out <= PPCMPLBWRDBUS_outdelay after OUT_DELAY;
	PPCS0PLBADDRACK_out <= PPCS0PLBADDRACK_outdelay after OUT_DELAY;
	PPCS0PLBMBUSY_out <= PPCS0PLBMBUSY_outdelay after OUT_DELAY;
	PPCS0PLBMIRQ_out <= PPCS0PLBMIRQ_outdelay after OUT_DELAY;
	PPCS0PLBMRDERR_out <= PPCS0PLBMRDERR_outdelay after OUT_DELAY;
	PPCS0PLBMWRERR_out <= PPCS0PLBMWRERR_outdelay after OUT_DELAY;
	PPCS0PLBRDBTERM_out <= PPCS0PLBRDBTERM_outdelay after OUT_DELAY;
	PPCS0PLBRDCOMP_out <= PPCS0PLBRDCOMP_outdelay after OUT_DELAY;
	PPCS0PLBRDDACK_out <= PPCS0PLBRDDACK_outdelay after OUT_DELAY;
	PPCS0PLBRDDBUS_out <= PPCS0PLBRDDBUS_outdelay after OUT_DELAY;
	PPCS0PLBRDWDADDR_out <= PPCS0PLBRDWDADDR_outdelay after OUT_DELAY;
	PPCS0PLBREARBITRATE_out <= PPCS0PLBREARBITRATE_outdelay after OUT_DELAY;
	PPCS0PLBSSIZE_out <= PPCS0PLBSSIZE_outdelay after OUT_DELAY;
	PPCS0PLBWAIT_out <= PPCS0PLBWAIT_outdelay after OUT_DELAY;
	PPCS0PLBWRBTERM_out <= PPCS0PLBWRBTERM_outdelay after OUT_DELAY;
	PPCS0PLBWRCOMP_out <= PPCS0PLBWRCOMP_outdelay after OUT_DELAY;
	PPCS0PLBWRDACK_out <= PPCS0PLBWRDACK_outdelay after OUT_DELAY;
	PPCS1PLBADDRACK_out <= PPCS1PLBADDRACK_outdelay after OUT_DELAY;
	PPCS1PLBMBUSY_out <= PPCS1PLBMBUSY_outdelay after OUT_DELAY;
	PPCS1PLBMIRQ_out <= PPCS1PLBMIRQ_outdelay after OUT_DELAY;
	PPCS1PLBMRDERR_out <= PPCS1PLBMRDERR_outdelay after OUT_DELAY;
	PPCS1PLBMWRERR_out <= PPCS1PLBMWRERR_outdelay after OUT_DELAY;
	PPCS1PLBRDBTERM_out <= PPCS1PLBRDBTERM_outdelay after OUT_DELAY;
	PPCS1PLBRDCOMP_out <= PPCS1PLBRDCOMP_outdelay after OUT_DELAY;
	PPCS1PLBRDDACK_out <= PPCS1PLBRDDACK_outdelay after OUT_DELAY;
	PPCS1PLBRDDBUS_out <= PPCS1PLBRDDBUS_outdelay after OUT_DELAY;
	PPCS1PLBRDWDADDR_out <= PPCS1PLBRDWDADDR_outdelay after OUT_DELAY;
	PPCS1PLBREARBITRATE_out <= PPCS1PLBREARBITRATE_outdelay after OUT_DELAY;
	PPCS1PLBSSIZE_out <= PPCS1PLBSSIZE_outdelay after OUT_DELAY;
	PPCS1PLBWAIT_out <= PPCS1PLBWAIT_outdelay after OUT_DELAY;
	PPCS1PLBWRBTERM_out <= PPCS1PLBWRBTERM_outdelay after OUT_DELAY;
	PPCS1PLBWRCOMP_out <= PPCS1PLBWRCOMP_outdelay after OUT_DELAY;
	PPCS1PLBWRDACK_out <= PPCS1PLBWRDACK_outdelay after OUT_DELAY;

	CPMC440CLK_indelay <= CPMC440CLK_dly after CLK_DELAY;
	CPMC440TIMERCLOCK_indelay <= CPMC440TIMERCLOCK_dly after CLK_DELAY;
	CPMDCRCLK_indelay <= CPMDCRCLK_dly after CLK_DELAY;
	CPMDMA0LLCLK_indelay <= CPMDMA0LLCLK_dly after CLK_DELAY;
	CPMDMA1LLCLK_indelay <= CPMDMA1LLCLK_dly after CLK_DELAY;
	CPMDMA2LLCLK_indelay <= CPMDMA2LLCLK_dly after CLK_DELAY;
	CPMDMA3LLCLK_indelay <= CPMDMA3LLCLK_dly after CLK_DELAY;
	CPMFCMCLK_indelay <= CPMFCMCLK_dly after CLK_DELAY;
	CPMINTERCONNECTCLK_indelay <= CPMINTERCONNECTCLK_dly after CLK_DELAY;
	CPMMCCLK_indelay <= CPMMCCLK_dly after CLK_DELAY;
	CPMPPCMPLBCLK_indelay <= CPMPPCMPLBCLK_dly after CLK_DELAY;
	CPMPPCS0PLBCLK_indelay <= CPMPPCS0PLBCLK_dly after CLK_DELAY;
	CPMPPCS1PLBCLK_indelay <= CPMPPCS1PLBCLK_dly after CLK_DELAY;
	JTGC440TCK_indelay <= JTGC440TCK_dly after CLK_DELAY;

	CPMC440CLKEN_indelay <= CPMC440CLKEN_dly after IN_DELAY;
	CPMC440CORECLOCKINACTIVE_indelay <= CPMC440CORECLOCKINACTIVE_dly after IN_DELAY;
	CPMINTERCONNECTCLKEN_indelay <= CPMINTERCONNECTCLKEN_dly after IN_DELAY;
	CPMINTERCONNECTCLKNTO1_indelay <= CPMINTERCONNECTCLKNTO1_dly after IN_DELAY;
	DBGC440DEBUGHALT_indelay <= DBGC440DEBUGHALT_dly after IN_DELAY;
	DBGC440SYSTEMSTATUS_indelay <= DBGC440SYSTEMSTATUS_dly after IN_DELAY;
	DBGC440UNCONDDEBUGEVENT_indelay <= DBGC440UNCONDDEBUGEVENT_dly after IN_DELAY;
	DCRPPCDMACK_indelay <= DCRPPCDMACK_dly after IN_DELAY;
	DCRPPCDMDBUSIN_indelay <= DCRPPCDMDBUSIN_dly after IN_DELAY;
	DCRPPCDMTIMEOUTWAIT_indelay <= DCRPPCDMTIMEOUTWAIT_dly after IN_DELAY;
	DCRPPCDSABUS_indelay <= DCRPPCDSABUS_dly after IN_DELAY;
	DCRPPCDSDBUSOUT_indelay <= DCRPPCDSDBUSOUT_dly after IN_DELAY;
	DCRPPCDSREAD_indelay <= DCRPPCDSREAD_dly after IN_DELAY;
	DCRPPCDSWRITE_indelay <= DCRPPCDSWRITE_dly after IN_DELAY;
	EICC440CRITIRQ_indelay <= EICC440CRITIRQ_dly after IN_DELAY;
	EICC440EXTIRQ_indelay <= EICC440EXTIRQ_dly after IN_DELAY;
	FCMAPUCONFIRMINSTR_indelay <= FCMAPUCONFIRMINSTR_dly after IN_DELAY;
	FCMAPUCR_indelay <= FCMAPUCR_dly after IN_DELAY;
	FCMAPUDONE_indelay <= FCMAPUDONE_dly after IN_DELAY;
	FCMAPUEXCEPTION_indelay <= FCMAPUEXCEPTION_dly after IN_DELAY;
	FCMAPUFPSCRFEX_indelay <= FCMAPUFPSCRFEX_dly after IN_DELAY;
	FCMAPURESULTVALID_indelay <= FCMAPURESULTVALID_dly after IN_DELAY;
	FCMAPURESULT_indelay <= FCMAPURESULT_dly after IN_DELAY;
	FCMAPUSLEEPNOTREADY_indelay <= FCMAPUSLEEPNOTREADY_dly after IN_DELAY;
	FCMAPUSTOREDATA_indelay <= FCMAPUSTOREDATA_dly after IN_DELAY;
	JTGC440TDI_indelay <= JTGC440TDI_dly after IN_DELAY;
	JTGC440TMS_indelay <= JTGC440TMS_dly after IN_DELAY;
	JTGC440TRSTNEG_indelay <= JTGC440TRSTNEG_dly after IN_DELAY;
	LLDMA0RSTENGINEREQ_indelay <= LLDMA0RSTENGINEREQ_dly after IN_DELAY;
	LLDMA0RXD_indelay <= LLDMA0RXD_dly after IN_DELAY;
	LLDMA0RXEOFN_indelay <= LLDMA0RXEOFN_dly after IN_DELAY;
	LLDMA0RXEOPN_indelay <= LLDMA0RXEOPN_dly after IN_DELAY;
	LLDMA0RXREM_indelay <= LLDMA0RXREM_dly after IN_DELAY;
	LLDMA0RXSOFN_indelay <= LLDMA0RXSOFN_dly after IN_DELAY;
	LLDMA0RXSOPN_indelay <= LLDMA0RXSOPN_dly after IN_DELAY;
	LLDMA0RXSRCRDYN_indelay <= LLDMA0RXSRCRDYN_dly after IN_DELAY;
	LLDMA0TXDSTRDYN_indelay <= LLDMA0TXDSTRDYN_dly after IN_DELAY;
	LLDMA1RSTENGINEREQ_indelay <= LLDMA1RSTENGINEREQ_dly after IN_DELAY;
	LLDMA1RXD_indelay <= LLDMA1RXD_dly after IN_DELAY;
	LLDMA1RXEOFN_indelay <= LLDMA1RXEOFN_dly after IN_DELAY;
	LLDMA1RXEOPN_indelay <= LLDMA1RXEOPN_dly after IN_DELAY;
	LLDMA1RXREM_indelay <= LLDMA1RXREM_dly after IN_DELAY;
	LLDMA1RXSOFN_indelay <= LLDMA1RXSOFN_dly after IN_DELAY;
	LLDMA1RXSOPN_indelay <= LLDMA1RXSOPN_dly after IN_DELAY;
	LLDMA1RXSRCRDYN_indelay <= LLDMA1RXSRCRDYN_dly after IN_DELAY;
	LLDMA1TXDSTRDYN_indelay <= LLDMA1TXDSTRDYN_dly after IN_DELAY;
	LLDMA2RSTENGINEREQ_indelay <= LLDMA2RSTENGINEREQ_dly after IN_DELAY;
	LLDMA2RXD_indelay <= LLDMA2RXD_dly after IN_DELAY;
	LLDMA2RXEOFN_indelay <= LLDMA2RXEOFN_dly after IN_DELAY;
	LLDMA2RXEOPN_indelay <= LLDMA2RXEOPN_dly after IN_DELAY;
	LLDMA2RXREM_indelay <= LLDMA2RXREM_dly after IN_DELAY;
	LLDMA2RXSOFN_indelay <= LLDMA2RXSOFN_dly after IN_DELAY;
	LLDMA2RXSOPN_indelay <= LLDMA2RXSOPN_dly after IN_DELAY;
	LLDMA2RXSRCRDYN_indelay <= LLDMA2RXSRCRDYN_dly after IN_DELAY;
	LLDMA2TXDSTRDYN_indelay <= LLDMA2TXDSTRDYN_dly after IN_DELAY;
	LLDMA3RSTENGINEREQ_indelay <= LLDMA3RSTENGINEREQ_dly after IN_DELAY;
	LLDMA3RXD_indelay <= LLDMA3RXD_dly after IN_DELAY;
	LLDMA3RXEOFN_indelay <= LLDMA3RXEOFN_dly after IN_DELAY;
	LLDMA3RXEOPN_indelay <= LLDMA3RXEOPN_dly after IN_DELAY;
	LLDMA3RXREM_indelay <= LLDMA3RXREM_dly after IN_DELAY;
	LLDMA3RXSOFN_indelay <= LLDMA3RXSOFN_dly after IN_DELAY;
	LLDMA3RXSOPN_indelay <= LLDMA3RXSOPN_dly after IN_DELAY;
	LLDMA3RXSRCRDYN_indelay <= LLDMA3RXSRCRDYN_dly after IN_DELAY;
	LLDMA3TXDSTRDYN_indelay <= LLDMA3TXDSTRDYN_dly after IN_DELAY;
	MCMIADDRREADYTOACCEPT_indelay <= MCMIADDRREADYTOACCEPT_dly after IN_DELAY;
	MCMIREADDATAERR_indelay <= MCMIREADDATAERR_dly after IN_DELAY;
	MCMIREADDATAVALID_indelay <= MCMIREADDATAVALID_dly after IN_DELAY;
	MCMIREADDATA_indelay <= MCMIREADDATA_dly after IN_DELAY;
	PLBPPCMADDRACK_indelay <= PLBPPCMADDRACK_dly after IN_DELAY;
	PLBPPCMMBUSY_indelay <= PLBPPCMMBUSY_dly after IN_DELAY;
	PLBPPCMMIRQ_indelay <= PLBPPCMMIRQ_dly after IN_DELAY;
	PLBPPCMMRDERR_indelay <= PLBPPCMMRDERR_dly after IN_DELAY;
	PLBPPCMMWRERR_indelay <= PLBPPCMMWRERR_dly after IN_DELAY;
	PLBPPCMRDBTERM_indelay <= PLBPPCMRDBTERM_dly after IN_DELAY;
	PLBPPCMRDDACK_indelay <= PLBPPCMRDDACK_dly after IN_DELAY;
	PLBPPCMRDDBUS_indelay <= PLBPPCMRDDBUS_dly after IN_DELAY;
	PLBPPCMRDPENDPRI_indelay <= PLBPPCMRDPENDPRI_dly after IN_DELAY;
	PLBPPCMRDPENDREQ_indelay <= PLBPPCMRDPENDREQ_dly after IN_DELAY;
	PLBPPCMRDWDADDR_indelay <= PLBPPCMRDWDADDR_dly after IN_DELAY;
	PLBPPCMREARBITRATE_indelay <= PLBPPCMREARBITRATE_dly after IN_DELAY;
	PLBPPCMREQPRI_indelay <= PLBPPCMREQPRI_dly after IN_DELAY;
	PLBPPCMSSIZE_indelay <= PLBPPCMSSIZE_dly after IN_DELAY;
	PLBPPCMTIMEOUT_indelay <= PLBPPCMTIMEOUT_dly after IN_DELAY;
	PLBPPCMWRBTERM_indelay <= PLBPPCMWRBTERM_dly after IN_DELAY;
	PLBPPCMWRDACK_indelay <= PLBPPCMWRDACK_dly after IN_DELAY;
	PLBPPCMWRPENDPRI_indelay <= PLBPPCMWRPENDPRI_dly after IN_DELAY;
	PLBPPCMWRPENDREQ_indelay <= PLBPPCMWRPENDREQ_dly after IN_DELAY;
	PLBPPCS0ABORT_indelay <= PLBPPCS0ABORT_dly after IN_DELAY;
	PLBPPCS0ABUS_indelay <= PLBPPCS0ABUS_dly after IN_DELAY;
	PLBPPCS0BE_indelay <= PLBPPCS0BE_dly after IN_DELAY;
	PLBPPCS0BUSLOCK_indelay <= PLBPPCS0BUSLOCK_dly after IN_DELAY;
	PLBPPCS0LOCKERR_indelay <= PLBPPCS0LOCKERR_dly after IN_DELAY;
	PLBPPCS0MASTERID_indelay <= PLBPPCS0MASTERID_dly after IN_DELAY;
	PLBPPCS0MSIZE_indelay <= PLBPPCS0MSIZE_dly after IN_DELAY;
	PLBPPCS0PAVALID_indelay <= PLBPPCS0PAVALID_dly after IN_DELAY;
	PLBPPCS0RDBURST_indelay <= PLBPPCS0RDBURST_dly after IN_DELAY;
	PLBPPCS0RDPENDPRI_indelay <= PLBPPCS0RDPENDPRI_dly after IN_DELAY;
	PLBPPCS0RDPENDREQ_indelay <= PLBPPCS0RDPENDREQ_dly after IN_DELAY;
	PLBPPCS0RDPRIM_indelay <= PLBPPCS0RDPRIM_dly after IN_DELAY;
	PLBPPCS0REQPRI_indelay <= PLBPPCS0REQPRI_dly after IN_DELAY;
	PLBPPCS0RNW_indelay <= PLBPPCS0RNW_dly after IN_DELAY;
	PLBPPCS0SAVALID_indelay <= PLBPPCS0SAVALID_dly after IN_DELAY;
	PLBPPCS0SIZE_indelay <= PLBPPCS0SIZE_dly after IN_DELAY;
	PLBPPCS0TATTRIBUTE_indelay <= PLBPPCS0TATTRIBUTE_dly after IN_DELAY;
	PLBPPCS0TYPE_indelay <= PLBPPCS0TYPE_dly after IN_DELAY;
	PLBPPCS0UABUS_indelay <= PLBPPCS0UABUS_dly after IN_DELAY;
	PLBPPCS0WRBURST_indelay <= PLBPPCS0WRBURST_dly after IN_DELAY;
	PLBPPCS0WRDBUS_indelay <= PLBPPCS0WRDBUS_dly after IN_DELAY;
	PLBPPCS0WRPENDPRI_indelay <= PLBPPCS0WRPENDPRI_dly after IN_DELAY;
	PLBPPCS0WRPENDREQ_indelay <= PLBPPCS0WRPENDREQ_dly after IN_DELAY;
	PLBPPCS0WRPRIM_indelay <= PLBPPCS0WRPRIM_dly after IN_DELAY;
	PLBPPCS1ABORT_indelay <= PLBPPCS1ABORT_dly after IN_DELAY;
	PLBPPCS1ABUS_indelay <= PLBPPCS1ABUS_dly after IN_DELAY;
	PLBPPCS1BE_indelay <= PLBPPCS1BE_dly after IN_DELAY;
	PLBPPCS1BUSLOCK_indelay <= PLBPPCS1BUSLOCK_dly after IN_DELAY;
	PLBPPCS1LOCKERR_indelay <= PLBPPCS1LOCKERR_dly after IN_DELAY;
	PLBPPCS1MASTERID_indelay <= PLBPPCS1MASTERID_dly after IN_DELAY;
	PLBPPCS1MSIZE_indelay <= PLBPPCS1MSIZE_dly after IN_DELAY;
	PLBPPCS1PAVALID_indelay <= PLBPPCS1PAVALID_dly after IN_DELAY;
	PLBPPCS1RDBURST_indelay <= PLBPPCS1RDBURST_dly after IN_DELAY;
	PLBPPCS1RDPENDPRI_indelay <= PLBPPCS1RDPENDPRI_dly after IN_DELAY;
	PLBPPCS1RDPENDREQ_indelay <= PLBPPCS1RDPENDREQ_dly after IN_DELAY;
	PLBPPCS1RDPRIM_indelay <= PLBPPCS1RDPRIM_dly after IN_DELAY;
	PLBPPCS1REQPRI_indelay <= PLBPPCS1REQPRI_dly after IN_DELAY;
	PLBPPCS1RNW_indelay <= PLBPPCS1RNW_dly after IN_DELAY;
	PLBPPCS1SAVALID_indelay <= PLBPPCS1SAVALID_dly after IN_DELAY;
	PLBPPCS1SIZE_indelay <= PLBPPCS1SIZE_dly after IN_DELAY;
	PLBPPCS1TATTRIBUTE_indelay <= PLBPPCS1TATTRIBUTE_dly after IN_DELAY;
	PLBPPCS1TYPE_indelay <= PLBPPCS1TYPE_dly after IN_DELAY;
	PLBPPCS1UABUS_indelay <= PLBPPCS1UABUS_dly after IN_DELAY;
	PLBPPCS1WRBURST_indelay <= PLBPPCS1WRBURST_dly after IN_DELAY;
	PLBPPCS1WRDBUS_indelay <= PLBPPCS1WRDBUS_dly after IN_DELAY;
	PLBPPCS1WRPENDPRI_indelay <= PLBPPCS1WRPENDPRI_dly after IN_DELAY;
	PLBPPCS1WRPENDREQ_indelay <= PLBPPCS1WRPENDREQ_dly after IN_DELAY;
	PLBPPCS1WRPRIM_indelay <= PLBPPCS1WRPRIM_dly after IN_DELAY;
	RSTC440RESETCHIP_indelay <= RSTC440RESETCHIP_dly after IN_DELAY;
	RSTC440RESETCORE_indelay <= RSTC440RESETCORE_dly after IN_DELAY;
	RSTC440RESETSYSTEM_indelay <= RSTC440RESETSYSTEM_dly after IN_DELAY;
	TIEC440DCURDLDCACHEPLBPRIO_indelay <= TIEC440DCURDLDCACHEPLBPRIO_dly after IN_DELAY;
	TIEC440DCURDNONCACHEPLBPRIO_indelay <= TIEC440DCURDNONCACHEPLBPRIO_dly after IN_DELAY;
	TIEC440DCURDTOUCHPLBPRIO_indelay <= TIEC440DCURDTOUCHPLBPRIO_dly after IN_DELAY;
	TIEC440DCURDURGENTPLBPRIO_indelay <= TIEC440DCURDURGENTPLBPRIO_dly after IN_DELAY;
	TIEC440DCUWRFLUSHPLBPRIO_indelay <= TIEC440DCUWRFLUSHPLBPRIO_dly after IN_DELAY;
	TIEC440DCUWRSTOREPLBPRIO_indelay <= TIEC440DCUWRSTOREPLBPRIO_dly after IN_DELAY;
	TIEC440DCUWRURGENTPLBPRIO_indelay <= TIEC440DCUWRURGENTPLBPRIO_dly after IN_DELAY;
	TIEC440ENDIANRESET_indelay <= TIEC440ENDIANRESET_dly after IN_DELAY;
	TIEC440ERPNRESET_indelay <= TIEC440ERPNRESET_dly after IN_DELAY;
	TIEC440ICURDFETCHPLBPRIO_indelay <= TIEC440ICURDFETCHPLBPRIO_dly after IN_DELAY;
	TIEC440ICURDSPECPLBPRIO_indelay <= TIEC440ICURDSPECPLBPRIO_dly after IN_DELAY;
	TIEC440ICURDTOUCHPLBPRIO_indelay <= TIEC440ICURDTOUCHPLBPRIO_dly after IN_DELAY;
	TIEC440PIR_indelay <= TIEC440PIR_dly after IN_DELAY;
	TIEC440PVR_indelay <= TIEC440PVR_dly after IN_DELAY;
	TIEC440USERRESET_indelay <= TIEC440USERRESET_dly after IN_DELAY;
	TIEDCRBASEADDR_indelay <= TIEDCRBASEADDR_dly after IN_DELAY;
	TRCC440TRACEDISABLE_indelay <= TRCC440TRACEDISABLE_dly after IN_DELAY;
	TRCC440TRIGGEREVENTIN_indelay <= TRCC440TRIGGEREVENTIN_dly after IN_DELAY;

	ppc440_swift_1 : PPC440_SWIFT
	port map (
	APU_CONTROL  =>  APU_CONTROL_BINARY,
	APU_UDI0  =>  APU_UDI0_BINARY,
	APU_UDI1  =>  APU_UDI1_BINARY,
	APU_UDI10  =>  APU_UDI10_BINARY,
	APU_UDI11  =>  APU_UDI11_BINARY,
	APU_UDI12  =>  APU_UDI12_BINARY,
	APU_UDI13  =>  APU_UDI13_BINARY,
	APU_UDI14  =>  APU_UDI14_BINARY,
	APU_UDI15  =>  APU_UDI15_BINARY,
	APU_UDI2  =>  APU_UDI2_BINARY,
	APU_UDI3  =>  APU_UDI3_BINARY,
	APU_UDI4  =>  APU_UDI4_BINARY,
	APU_UDI5  =>  APU_UDI5_BINARY,
	APU_UDI6  =>  APU_UDI6_BINARY,
	APU_UDI7  =>  APU_UDI7_BINARY,
	APU_UDI8  =>  APU_UDI8_BINARY,
	APU_UDI9  =>  APU_UDI9_BINARY,
	CLOCK_DELAY  =>  CLOCK_DELAY_BINARY,
	DCR_AUTOLOCK_ENABLE  =>  DCR_AUTOLOCK_ENABLE_BINARY,
	DMA0_CONTROL  =>  DMA0_CONTROL_BINARY,
	DMA0_RXCHANNELCTRL  =>  DMA0_RXCHANNELCTRL_BINARY,
	DMA0_RXIRQTIMER  =>  DMA0_RXIRQTIMER_BINARY,
	DMA0_TXCHANNELCTRL  =>  DMA0_TXCHANNELCTRL_BINARY,
	DMA0_TXIRQTIMER  =>  DMA0_TXIRQTIMER_BINARY,
	DMA1_CONTROL  =>  DMA1_CONTROL_BINARY,
	DMA1_RXCHANNELCTRL  =>  DMA1_RXCHANNELCTRL_BINARY,
	DMA1_RXIRQTIMER  =>  DMA1_RXIRQTIMER_BINARY,
	DMA1_TXCHANNELCTRL  =>  DMA1_TXCHANNELCTRL_BINARY,
	DMA1_TXIRQTIMER  =>  DMA1_TXIRQTIMER_BINARY,
	DMA2_CONTROL  =>  DMA2_CONTROL_BINARY,
	DMA2_RXCHANNELCTRL  =>  DMA2_RXCHANNELCTRL_BINARY,
	DMA2_RXIRQTIMER  =>  DMA2_RXIRQTIMER_BINARY,
	DMA2_TXCHANNELCTRL  =>  DMA2_TXCHANNELCTRL_BINARY,
	DMA2_TXIRQTIMER  =>  DMA2_TXIRQTIMER_BINARY,
	DMA3_CONTROL  =>  DMA3_CONTROL_BINARY,
	DMA3_RXCHANNELCTRL  =>  DMA3_RXCHANNELCTRL_BINARY,
	DMA3_RXIRQTIMER  =>  DMA3_RXIRQTIMER_BINARY,
	DMA3_TXCHANNELCTRL  =>  DMA3_TXCHANNELCTRL_BINARY,
	DMA3_TXIRQTIMER  =>  DMA3_TXIRQTIMER_BINARY,
	INTERCONNECT_IMASK  =>  INTERCONNECT_IMASK_BINARY,
	INTERCONNECT_TMPL_SEL  =>  INTERCONNECT_TMPL_SEL_BINARY,
	MI_ARBCONFIG  =>  MI_ARBCONFIG_BINARY,
	MI_BANKCONFLICT_MASK  =>  MI_BANKCONFLICT_MASK_BINARY,
	MI_CONTROL  =>  MI_CONTROL_BINARY,
	MI_ROWCONFLICT_MASK  =>  MI_ROWCONFLICT_MASK_BINARY,
	PPCDM_ASYNCMODE  =>  PPCDM_ASYNCMODE_BINARY,
	PPCDS_ASYNCMODE  =>  PPCDS_ASYNCMODE_BINARY,
	PPCM_ARBCONFIG  =>  PPCM_ARBCONFIG_BINARY,
	PPCM_CONTROL  =>  PPCM_CONTROL_BINARY,
	PPCM_COUNTER  =>  PPCM_COUNTER_BINARY,
	PPCS0_ADDRMAP_TMPL0  =>  PPCS0_ADDRMAP_TMPL0_BINARY,
	PPCS0_ADDRMAP_TMPL1  =>  PPCS0_ADDRMAP_TMPL1_BINARY,
	PPCS0_ADDRMAP_TMPL2  =>  PPCS0_ADDRMAP_TMPL2_BINARY,
	PPCS0_ADDRMAP_TMPL3  =>  PPCS0_ADDRMAP_TMPL3_BINARY,
	PPCS0_CONTROL  =>  PPCS0_CONTROL_BINARY,
	PPCS0_WIDTH_128N64  =>  PPCS0_WIDTH_128N64_BINARY,
	PPCS1_ADDRMAP_TMPL0  =>  PPCS1_ADDRMAP_TMPL0_BINARY,
	PPCS1_ADDRMAP_TMPL1  =>  PPCS1_ADDRMAP_TMPL1_BINARY,
	PPCS1_ADDRMAP_TMPL2  =>  PPCS1_ADDRMAP_TMPL2_BINARY,
	PPCS1_ADDRMAP_TMPL3  =>  PPCS1_ADDRMAP_TMPL3_BINARY,
	PPCS1_CONTROL  =>  PPCS1_CONTROL_BINARY,
	PPCS1_WIDTH_128N64  =>  PPCS1_WIDTH_128N64_BINARY,
	XBAR_ADDRMAP_TMPL0  =>  XBAR_ADDRMAP_TMPL0_BINARY,
	XBAR_ADDRMAP_TMPL1  =>  XBAR_ADDRMAP_TMPL1_BINARY,
	XBAR_ADDRMAP_TMPL2  =>  XBAR_ADDRMAP_TMPL2_BINARY,
	XBAR_ADDRMAP_TMPL3  =>  XBAR_ADDRMAP_TMPL3_BINARY,

	APUFCMDECFPUOP  =>  APUFCMDECFPUOP_outdelay,
	APUFCMDECLDSTXFERSIZE  =>  APUFCMDECLDSTXFERSIZE_outdelay,
	APUFCMDECLOAD  =>  APUFCMDECLOAD_outdelay,
	APUFCMDECNONAUTON  =>  APUFCMDECNONAUTON_outdelay,
	APUFCMDECSTORE  =>  APUFCMDECSTORE_outdelay,
	APUFCMDECUDI  =>  APUFCMDECUDI_outdelay,
	APUFCMDECUDIVALID  =>  APUFCMDECUDIVALID_outdelay,
	APUFCMENDIAN  =>  APUFCMENDIAN_outdelay,
	APUFCMFLUSH  =>  APUFCMFLUSH_outdelay,
	APUFCMINSTRUCTION  =>  APUFCMINSTRUCTION_outdelay,
	APUFCMINSTRVALID  =>  APUFCMINSTRVALID_outdelay,
	APUFCMLOADBYTEADDR  =>  APUFCMLOADBYTEADDR_outdelay,
	APUFCMLOADDATA  =>  APUFCMLOADDATA_outdelay,
	APUFCMLOADDVALID  =>  APUFCMLOADDVALID_outdelay,
	APUFCMMSRFE0  =>  APUFCMMSRFE0_outdelay,
	APUFCMMSRFE1  =>  APUFCMMSRFE1_outdelay,
	APUFCMNEXTINSTRREADY  =>  APUFCMNEXTINSTRREADY_outdelay,
	APUFCMOPERANDVALID  =>  APUFCMOPERANDVALID_outdelay,
	APUFCMRADATA  =>  APUFCMRADATA_outdelay,
	APUFCMRBDATA  =>  APUFCMRBDATA_outdelay,
	APUFCMWRITEBACKOK  =>  APUFCMWRITEBACKOK_outdelay,
	C440CPMCORESLEEPREQ  =>  C440CPMCORESLEEPREQ_outdelay,
	C440CPMDECIRPTREQ  =>  C440CPMDECIRPTREQ_outdelay,
	C440CPMFITIRPTREQ  =>  C440CPMFITIRPTREQ_outdelay,
	C440CPMMSRCE  =>  C440CPMMSRCE_outdelay,
	C440CPMMSREE  =>  C440CPMMSREE_outdelay,
	C440CPMTIMERRESETREQ  =>  C440CPMTIMERRESETREQ_outdelay,
	C440CPMWDIRPTREQ  =>  C440CPMWDIRPTREQ_outdelay,
	C440DBGSYSTEMCONTROL  =>  C440DBGSYSTEMCONTROL_outdelay,
	C440JTGTDO  =>  C440JTGTDO_outdelay,
	C440JTGTDOEN  =>  C440JTGTDOEN_outdelay,
	C440MACHINECHECK  =>  C440MACHINECHECK_outdelay,
	C440RSTCHIPRESETREQ  =>  C440RSTCHIPRESETREQ_outdelay,
	C440RSTCORERESETREQ  =>  C440RSTCORERESETREQ_outdelay,
	C440RSTSYSTEMRESETREQ  =>  C440RSTSYSTEMRESETREQ_outdelay,
	C440TRCBRANCHSTATUS  =>  C440TRCBRANCHSTATUS_outdelay,
	C440TRCCYCLE  =>  C440TRCCYCLE_outdelay,
	C440TRCEXECUTIONSTATUS  =>  C440TRCEXECUTIONSTATUS_outdelay,
	C440TRCTRACESTATUS  =>  C440TRCTRACESTATUS_outdelay,
	C440TRCTRIGGEREVENTOUT  =>  C440TRCTRIGGEREVENTOUT_outdelay,
	C440TRCTRIGGEREVENTTYPE  =>  C440TRCTRIGGEREVENTTYPE_outdelay,
	DMA0LLRSTENGINEACK  =>  DMA0LLRSTENGINEACK_outdelay,
	DMA0LLRXDSTRDYN  =>  DMA0LLRXDSTRDYN_outdelay,
	DMA0LLTXD  =>  DMA0LLTXD_outdelay,
	DMA0LLTXEOFN  =>  DMA0LLTXEOFN_outdelay,
	DMA0LLTXEOPN  =>  DMA0LLTXEOPN_outdelay,
	DMA0LLTXREM  =>  DMA0LLTXREM_outdelay,
	DMA0LLTXSOFN  =>  DMA0LLTXSOFN_outdelay,
	DMA0LLTXSOPN  =>  DMA0LLTXSOPN_outdelay,
	DMA0LLTXSRCRDYN  =>  DMA0LLTXSRCRDYN_outdelay,
	DMA0RXIRQ  =>  DMA0RXIRQ_outdelay,
	DMA0TXIRQ  =>  DMA0TXIRQ_outdelay,
	DMA1LLRSTENGINEACK  =>  DMA1LLRSTENGINEACK_outdelay,
	DMA1LLRXDSTRDYN  =>  DMA1LLRXDSTRDYN_outdelay,
	DMA1LLTXD  =>  DMA1LLTXD_outdelay,
	DMA1LLTXEOFN  =>  DMA1LLTXEOFN_outdelay,
	DMA1LLTXEOPN  =>  DMA1LLTXEOPN_outdelay,
	DMA1LLTXREM  =>  DMA1LLTXREM_outdelay,
	DMA1LLTXSOFN  =>  DMA1LLTXSOFN_outdelay,
	DMA1LLTXSOPN  =>  DMA1LLTXSOPN_outdelay,
	DMA1LLTXSRCRDYN  =>  DMA1LLTXSRCRDYN_outdelay,
	DMA1RXIRQ  =>  DMA1RXIRQ_outdelay,
	DMA1TXIRQ  =>  DMA1TXIRQ_outdelay,
	DMA2LLRSTENGINEACK  =>  DMA2LLRSTENGINEACK_outdelay,
	DMA2LLRXDSTRDYN  =>  DMA2LLRXDSTRDYN_outdelay,
	DMA2LLTXD  =>  DMA2LLTXD_outdelay,
	DMA2LLTXEOFN  =>  DMA2LLTXEOFN_outdelay,
	DMA2LLTXEOPN  =>  DMA2LLTXEOPN_outdelay,
	DMA2LLTXREM  =>  DMA2LLTXREM_outdelay,
	DMA2LLTXSOFN  =>  DMA2LLTXSOFN_outdelay,
	DMA2LLTXSOPN  =>  DMA2LLTXSOPN_outdelay,
	DMA2LLTXSRCRDYN  =>  DMA2LLTXSRCRDYN_outdelay,
	DMA2RXIRQ  =>  DMA2RXIRQ_outdelay,
	DMA2TXIRQ  =>  DMA2TXIRQ_outdelay,
	DMA3LLRSTENGINEACK  =>  DMA3LLRSTENGINEACK_outdelay,
	DMA3LLRXDSTRDYN  =>  DMA3LLRXDSTRDYN_outdelay,
	DMA3LLTXD  =>  DMA3LLTXD_outdelay,
	DMA3LLTXEOFN  =>  DMA3LLTXEOFN_outdelay,
	DMA3LLTXEOPN  =>  DMA3LLTXEOPN_outdelay,
	DMA3LLTXREM  =>  DMA3LLTXREM_outdelay,
	DMA3LLTXSOFN  =>  DMA3LLTXSOFN_outdelay,
	DMA3LLTXSOPN  =>  DMA3LLTXSOPN_outdelay,
	DMA3LLTXSRCRDYN  =>  DMA3LLTXSRCRDYN_outdelay,
	DMA3RXIRQ  =>  DMA3RXIRQ_outdelay,
	DMA3TXIRQ  =>  DMA3TXIRQ_outdelay,
	MIMCADDRESS  =>  MIMCADDRESS_outdelay,
	MIMCADDRESSVALID  =>  MIMCADDRESSVALID_outdelay,
	MIMCBANKCONFLICT  =>  MIMCBANKCONFLICT_outdelay,
	MIMCBYTEENABLE  =>  MIMCBYTEENABLE_outdelay,
	MIMCREADNOTWRITE  =>  MIMCREADNOTWRITE_outdelay,
	MIMCROWCONFLICT  =>  MIMCROWCONFLICT_outdelay,
	MIMCWRITEDATA  =>  MIMCWRITEDATA_outdelay,
	MIMCWRITEDATAVALID  =>  MIMCWRITEDATAVALID_outdelay,
	PPCCPMINTERCONNECTBUSY  =>  PPCCPMINTERCONNECTBUSY_outdelay,
	PPCDMDCRABUS  =>  PPCDMDCRABUS_outdelay,
	PPCDMDCRDBUSOUT  =>  PPCDMDCRDBUSOUT_outdelay,
	PPCDMDCRREAD  =>  PPCDMDCRREAD_outdelay,
	PPCDMDCRUABUS  =>  PPCDMDCRUABUS_outdelay,
	PPCDMDCRWRITE  =>  PPCDMDCRWRITE_outdelay,
	PPCDSDCRACK  =>  PPCDSDCRACK_outdelay,
	PPCDSDCRDBUSIN  =>  PPCDSDCRDBUSIN_outdelay,
	PPCDSDCRTIMEOUTWAIT  =>  PPCDSDCRTIMEOUTWAIT_outdelay,
	PPCEICINTERCONNECTIRQ  =>  PPCEICINTERCONNECTIRQ_outdelay,
	PPCMPLBABORT  =>  PPCMPLBABORT_outdelay,
	PPCMPLBABUS  =>  PPCMPLBABUS_outdelay,
	PPCMPLBBE  =>  PPCMPLBBE_outdelay,
	PPCMPLBBUSLOCK  =>  PPCMPLBBUSLOCK_outdelay,
	PPCMPLBLOCKERR  =>  PPCMPLBLOCKERR_outdelay,
	PPCMPLBPRIORITY  =>  PPCMPLBPRIORITY_outdelay,
	PPCMPLBRDBURST  =>  PPCMPLBRDBURST_outdelay,
	PPCMPLBREQUEST  =>  PPCMPLBREQUEST_outdelay,
	PPCMPLBRNW  =>  PPCMPLBRNW_outdelay,
	PPCMPLBSIZE  =>  PPCMPLBSIZE_outdelay,
	PPCMPLBTATTRIBUTE  =>  PPCMPLBTATTRIBUTE_outdelay,
	PPCMPLBTYPE  =>  PPCMPLBTYPE_outdelay,
	PPCMPLBUABUS  =>  PPCMPLBUABUS_outdelay,
	PPCMPLBWRBURST  =>  PPCMPLBWRBURST_outdelay,
	PPCMPLBWRDBUS  =>  PPCMPLBWRDBUS_outdelay,
	PPCS0PLBADDRACK  =>  PPCS0PLBADDRACK_outdelay,
	PPCS0PLBMBUSY  =>  PPCS0PLBMBUSY_outdelay,
	PPCS0PLBMIRQ  =>  PPCS0PLBMIRQ_outdelay,
	PPCS0PLBMRDERR  =>  PPCS0PLBMRDERR_outdelay,
	PPCS0PLBMWRERR  =>  PPCS0PLBMWRERR_outdelay,
	PPCS0PLBRDBTERM  =>  PPCS0PLBRDBTERM_outdelay,
	PPCS0PLBRDCOMP  =>  PPCS0PLBRDCOMP_outdelay,
	PPCS0PLBRDDACK  =>  PPCS0PLBRDDACK_outdelay,
	PPCS0PLBRDDBUS  =>  PPCS0PLBRDDBUS_outdelay,
	PPCS0PLBRDWDADDR  =>  PPCS0PLBRDWDADDR_outdelay,
	PPCS0PLBREARBITRATE  =>  PPCS0PLBREARBITRATE_outdelay,
	PPCS0PLBSSIZE  =>  PPCS0PLBSSIZE_outdelay,
	PPCS0PLBWAIT  =>  PPCS0PLBWAIT_outdelay,
	PPCS0PLBWRBTERM  =>  PPCS0PLBWRBTERM_outdelay,
	PPCS0PLBWRCOMP  =>  PPCS0PLBWRCOMP_outdelay,
	PPCS0PLBWRDACK  =>  PPCS0PLBWRDACK_outdelay,
	PPCS1PLBADDRACK  =>  PPCS1PLBADDRACK_outdelay,
	PPCS1PLBMBUSY  =>  PPCS1PLBMBUSY_outdelay,
	PPCS1PLBMIRQ  =>  PPCS1PLBMIRQ_outdelay,
	PPCS1PLBMRDERR  =>  PPCS1PLBMRDERR_outdelay,
	PPCS1PLBMWRERR  =>  PPCS1PLBMWRERR_outdelay,
	PPCS1PLBRDBTERM  =>  PPCS1PLBRDBTERM_outdelay,
	PPCS1PLBRDCOMP  =>  PPCS1PLBRDCOMP_outdelay,
	PPCS1PLBRDDACK  =>  PPCS1PLBRDDACK_outdelay,
	PPCS1PLBRDDBUS  =>  PPCS1PLBRDDBUS_outdelay,
	PPCS1PLBRDWDADDR  =>  PPCS1PLBRDWDADDR_outdelay,
	PPCS1PLBREARBITRATE  =>  PPCS1PLBREARBITRATE_outdelay,
	PPCS1PLBSSIZE  =>  PPCS1PLBSSIZE_outdelay,
	PPCS1PLBWAIT  =>  PPCS1PLBWAIT_outdelay,
	PPCS1PLBWRBTERM  =>  PPCS1PLBWRBTERM_outdelay,
	PPCS1PLBWRCOMP  =>  PPCS1PLBWRCOMP_outdelay,
	PPCS1PLBWRDACK  =>  PPCS1PLBWRDACK_outdelay,

	CPMC440CLK  =>  CPMC440CLK_indelay,
	CPMC440CLKEN  =>  CPMC440CLKEN_indelay,
	CPMC440CORECLOCKINACTIVE  =>  CPMC440CORECLOCKINACTIVE_indelay,
	CPMC440TIMERCLOCK  =>  CPMC440TIMERCLOCK_indelay,
	CPMDCRCLK  =>  CPMDCRCLK_indelay,
	CPMDMA0LLCLK  =>  CPMDMA0LLCLK_indelay,
	CPMDMA1LLCLK  =>  CPMDMA1LLCLK_indelay,
	CPMDMA2LLCLK  =>  CPMDMA2LLCLK_indelay,
	CPMDMA3LLCLK  =>  CPMDMA3LLCLK_indelay,
	CPMFCMCLK  =>  CPMFCMCLK_indelay,
	CPMINTERCONNECTCLK  =>  CPMINTERCONNECTCLK_indelay,
	CPMINTERCONNECTCLKEN  =>  CPMINTERCONNECTCLKEN_indelay,
	CPMINTERCONNECTCLKNTO1  =>  CPMINTERCONNECTCLKNTO1_indelay,
	CPMMCCLK  =>  CPMMCCLK_indelay,
	CPMPPCMPLBCLK  =>  CPMPPCMPLBCLK_indelay,
	CPMPPCS0PLBCLK  =>  CPMPPCS0PLBCLK_indelay,
	CPMPPCS1PLBCLK  =>  CPMPPCS1PLBCLK_indelay,
	DBGC440DEBUGHALT  =>  DBGC440DEBUGHALT_indelay,
	DBGC440SYSTEMSTATUS  =>  DBGC440SYSTEMSTATUS_indelay,
	DBGC440UNCONDDEBUGEVENT  =>  DBGC440UNCONDDEBUGEVENT_indelay,
	DCRPPCDMACK  =>  DCRPPCDMACK_indelay,
	DCRPPCDMDBUSIN  =>  DCRPPCDMDBUSIN_indelay,
	DCRPPCDMTIMEOUTWAIT  =>  DCRPPCDMTIMEOUTWAIT_indelay,
	DCRPPCDSABUS  =>  DCRPPCDSABUS_indelay,
	DCRPPCDSDBUSOUT  =>  DCRPPCDSDBUSOUT_indelay,
	DCRPPCDSREAD  =>  DCRPPCDSREAD_indelay,
	DCRPPCDSWRITE  =>  DCRPPCDSWRITE_indelay,
	EICC440CRITIRQ  =>  EICC440CRITIRQ_indelay,
	EICC440EXTIRQ  =>  EICC440EXTIRQ_indelay,
	FCMAPUCONFIRMINSTR  =>  FCMAPUCONFIRMINSTR_indelay,
	FCMAPUCR  =>  FCMAPUCR_indelay,
	FCMAPUDONE  =>  FCMAPUDONE_indelay,
	FCMAPUEXCEPTION  =>  FCMAPUEXCEPTION_indelay,
	FCMAPUFPSCRFEX  =>  FCMAPUFPSCRFEX_indelay,
	FCMAPURESULT  =>  FCMAPURESULT_indelay,
	FCMAPURESULTVALID  =>  FCMAPURESULTVALID_indelay,
	FCMAPUSLEEPNOTREADY  =>  FCMAPUSLEEPNOTREADY_indelay,
	FCMAPUSTOREDATA  =>  FCMAPUSTOREDATA_indelay,
	GSR  =>  GSR,
	JTGC440TCK  =>  JTGC440TCK_indelay,
	JTGC440TDI  =>  JTGC440TDI_indelay,
	JTGC440TMS  =>  JTGC440TMS_indelay,
	JTGC440TRSTNEG  =>  JTGC440TRSTNEG_indelay,
	LLDMA0RSTENGINEREQ  =>  LLDMA0RSTENGINEREQ_indelay,
	LLDMA0RXD  =>  LLDMA0RXD_indelay,
	LLDMA0RXEOFN  =>  LLDMA0RXEOFN_indelay,
	LLDMA0RXEOPN  =>  LLDMA0RXEOPN_indelay,
	LLDMA0RXREM  =>  LLDMA0RXREM_indelay,
	LLDMA0RXSOFN  =>  LLDMA0RXSOFN_indelay,
	LLDMA0RXSOPN  =>  LLDMA0RXSOPN_indelay,
	LLDMA0RXSRCRDYN  =>  LLDMA0RXSRCRDYN_indelay,
	LLDMA0TXDSTRDYN  =>  LLDMA0TXDSTRDYN_indelay,
	LLDMA1RSTENGINEREQ  =>  LLDMA1RSTENGINEREQ_indelay,
	LLDMA1RXD  =>  LLDMA1RXD_indelay,
	LLDMA1RXEOFN  =>  LLDMA1RXEOFN_indelay,
	LLDMA1RXEOPN  =>  LLDMA1RXEOPN_indelay,
	LLDMA1RXREM  =>  LLDMA1RXREM_indelay,
	LLDMA1RXSOFN  =>  LLDMA1RXSOFN_indelay,
	LLDMA1RXSOPN  =>  LLDMA1RXSOPN_indelay,
	LLDMA1RXSRCRDYN  =>  LLDMA1RXSRCRDYN_indelay,
	LLDMA1TXDSTRDYN  =>  LLDMA1TXDSTRDYN_indelay,
	LLDMA2RSTENGINEREQ  =>  LLDMA2RSTENGINEREQ_indelay,
	LLDMA2RXD  =>  LLDMA2RXD_indelay,
	LLDMA2RXEOFN  =>  LLDMA2RXEOFN_indelay,
	LLDMA2RXEOPN  =>  LLDMA2RXEOPN_indelay,
	LLDMA2RXREM  =>  LLDMA2RXREM_indelay,
	LLDMA2RXSOFN  =>  LLDMA2RXSOFN_indelay,
	LLDMA2RXSOPN  =>  LLDMA2RXSOPN_indelay,
	LLDMA2RXSRCRDYN  =>  LLDMA2RXSRCRDYN_indelay,
	LLDMA2TXDSTRDYN  =>  LLDMA2TXDSTRDYN_indelay,
	LLDMA3RSTENGINEREQ  =>  LLDMA3RSTENGINEREQ_indelay,
	LLDMA3RXD  =>  LLDMA3RXD_indelay,
	LLDMA3RXEOFN  =>  LLDMA3RXEOFN_indelay,
	LLDMA3RXEOPN  =>  LLDMA3RXEOPN_indelay,
	LLDMA3RXREM  =>  LLDMA3RXREM_indelay,
	LLDMA3RXSOFN  =>  LLDMA3RXSOFN_indelay,
	LLDMA3RXSOPN  =>  LLDMA3RXSOPN_indelay,
	LLDMA3RXSRCRDYN  =>  LLDMA3RXSRCRDYN_indelay,
	LLDMA3TXDSTRDYN  =>  LLDMA3TXDSTRDYN_indelay,
	MCMIADDRREADYTOACCEPT  =>  MCMIADDRREADYTOACCEPT_indelay,
	MCMIREADDATA  =>  MCMIREADDATA_indelay,
	MCMIREADDATAERR  =>  MCMIREADDATAERR_indelay,
	MCMIREADDATAVALID  =>  MCMIREADDATAVALID_indelay,
	PLBPPCMADDRACK  =>  PLBPPCMADDRACK_indelay,
	PLBPPCMMBUSY  =>  PLBPPCMMBUSY_indelay,
	PLBPPCMMIRQ  =>  PLBPPCMMIRQ_indelay,
	PLBPPCMMRDERR  =>  PLBPPCMMRDERR_indelay,
	PLBPPCMMWRERR  =>  PLBPPCMMWRERR_indelay,
	PLBPPCMRDBTERM  =>  PLBPPCMRDBTERM_indelay,
	PLBPPCMRDDACK  =>  PLBPPCMRDDACK_indelay,
	PLBPPCMRDDBUS  =>  PLBPPCMRDDBUS_indelay,
	PLBPPCMRDPENDPRI  =>  PLBPPCMRDPENDPRI_indelay,
	PLBPPCMRDPENDREQ  =>  PLBPPCMRDPENDREQ_indelay,
	PLBPPCMRDWDADDR  =>  PLBPPCMRDWDADDR_indelay,
	PLBPPCMREARBITRATE  =>  PLBPPCMREARBITRATE_indelay,
	PLBPPCMREQPRI  =>  PLBPPCMREQPRI_indelay,
	PLBPPCMSSIZE  =>  PLBPPCMSSIZE_indelay,
	PLBPPCMTIMEOUT  =>  PLBPPCMTIMEOUT_indelay,
	PLBPPCMWRBTERM  =>  PLBPPCMWRBTERM_indelay,
	PLBPPCMWRDACK  =>  PLBPPCMWRDACK_indelay,
	PLBPPCMWRPENDPRI  =>  PLBPPCMWRPENDPRI_indelay,
	PLBPPCMWRPENDREQ  =>  PLBPPCMWRPENDREQ_indelay,
	PLBPPCS0ABORT  =>  PLBPPCS0ABORT_indelay,
	PLBPPCS0ABUS  =>  PLBPPCS0ABUS_indelay,
	PLBPPCS0BE  =>  PLBPPCS0BE_indelay,
	PLBPPCS0BUSLOCK  =>  PLBPPCS0BUSLOCK_indelay,
	PLBPPCS0LOCKERR  =>  PLBPPCS0LOCKERR_indelay,
	PLBPPCS0MASTERID  =>  PLBPPCS0MASTERID_indelay,
	PLBPPCS0MSIZE  =>  PLBPPCS0MSIZE_indelay,
	PLBPPCS0PAVALID  =>  PLBPPCS0PAVALID_indelay,
	PLBPPCS0RDBURST  =>  PLBPPCS0RDBURST_indelay,
	PLBPPCS0RDPENDPRI  =>  PLBPPCS0RDPENDPRI_indelay,
	PLBPPCS0RDPENDREQ  =>  PLBPPCS0RDPENDREQ_indelay,
	PLBPPCS0RDPRIM  =>  PLBPPCS0RDPRIM_indelay,
	PLBPPCS0REQPRI  =>  PLBPPCS0REQPRI_indelay,
	PLBPPCS0RNW  =>  PLBPPCS0RNW_indelay,
	PLBPPCS0SAVALID  =>  PLBPPCS0SAVALID_indelay,
	PLBPPCS0SIZE  =>  PLBPPCS0SIZE_indelay,
	PLBPPCS0TATTRIBUTE  =>  PLBPPCS0TATTRIBUTE_indelay,
	PLBPPCS0TYPE  =>  PLBPPCS0TYPE_indelay,
	PLBPPCS0UABUS  =>  PLBPPCS0UABUS_indelay,
	PLBPPCS0WRBURST  =>  PLBPPCS0WRBURST_indelay,
	PLBPPCS0WRDBUS  =>  PLBPPCS0WRDBUS_indelay,
	PLBPPCS0WRPENDPRI  =>  PLBPPCS0WRPENDPRI_indelay,
	PLBPPCS0WRPENDREQ  =>  PLBPPCS0WRPENDREQ_indelay,
	PLBPPCS0WRPRIM  =>  PLBPPCS0WRPRIM_indelay,
	PLBPPCS1ABORT  =>  PLBPPCS1ABORT_indelay,
	PLBPPCS1ABUS  =>  PLBPPCS1ABUS_indelay,
	PLBPPCS1BE  =>  PLBPPCS1BE_indelay,
	PLBPPCS1BUSLOCK  =>  PLBPPCS1BUSLOCK_indelay,
	PLBPPCS1LOCKERR  =>  PLBPPCS1LOCKERR_indelay,
	PLBPPCS1MASTERID  =>  PLBPPCS1MASTERID_indelay,
	PLBPPCS1MSIZE  =>  PLBPPCS1MSIZE_indelay,
	PLBPPCS1PAVALID  =>  PLBPPCS1PAVALID_indelay,
	PLBPPCS1RDBURST  =>  PLBPPCS1RDBURST_indelay,
	PLBPPCS1RDPENDPRI  =>  PLBPPCS1RDPENDPRI_indelay,
	PLBPPCS1RDPENDREQ  =>  PLBPPCS1RDPENDREQ_indelay,
	PLBPPCS1RDPRIM  =>  PLBPPCS1RDPRIM_indelay,
	PLBPPCS1REQPRI  =>  PLBPPCS1REQPRI_indelay,
	PLBPPCS1RNW  =>  PLBPPCS1RNW_indelay,
	PLBPPCS1SAVALID  =>  PLBPPCS1SAVALID_indelay,
	PLBPPCS1SIZE  =>  PLBPPCS1SIZE_indelay,
	PLBPPCS1TATTRIBUTE  =>  PLBPPCS1TATTRIBUTE_indelay,
	PLBPPCS1TYPE  =>  PLBPPCS1TYPE_indelay,
	PLBPPCS1UABUS  =>  PLBPPCS1UABUS_indelay,
	PLBPPCS1WRBURST  =>  PLBPPCS1WRBURST_indelay,
	PLBPPCS1WRDBUS  =>  PLBPPCS1WRDBUS_indelay,
	PLBPPCS1WRPENDPRI  =>  PLBPPCS1WRPENDPRI_indelay,
	PLBPPCS1WRPENDREQ  =>  PLBPPCS1WRPENDREQ_indelay,
	PLBPPCS1WRPRIM  =>  PLBPPCS1WRPRIM_indelay,
	RSTC440RESETCHIP  =>  RSTC440RESETCHIP_indelay,
	RSTC440RESETCORE  =>  RSTC440RESETCORE_indelay,
	RSTC440RESETSYSTEM  =>  RSTC440RESETSYSTEM_indelay,
	TIEC440DCURDLDCACHEPLBPRIO  =>  TIEC440DCURDLDCACHEPLBPRIO_indelay,
	TIEC440DCURDNONCACHEPLBPRIO  =>  TIEC440DCURDNONCACHEPLBPRIO_indelay,
	TIEC440DCURDTOUCHPLBPRIO  =>  TIEC440DCURDTOUCHPLBPRIO_indelay,
	TIEC440DCURDURGENTPLBPRIO  =>  TIEC440DCURDURGENTPLBPRIO_indelay,
	TIEC440DCUWRFLUSHPLBPRIO  =>  TIEC440DCUWRFLUSHPLBPRIO_indelay,
	TIEC440DCUWRSTOREPLBPRIO  =>  TIEC440DCUWRSTOREPLBPRIO_indelay,
	TIEC440DCUWRURGENTPLBPRIO  =>  TIEC440DCUWRURGENTPLBPRIO_indelay,
	TIEC440ENDIANRESET  =>  TIEC440ENDIANRESET_indelay,
	TIEC440ERPNRESET  =>  TIEC440ERPNRESET_indelay,
	TIEC440ICURDFETCHPLBPRIO  =>  TIEC440ICURDFETCHPLBPRIO_indelay,
	TIEC440ICURDSPECPLBPRIO  =>  TIEC440ICURDSPECPLBPRIO_indelay,
	TIEC440ICURDTOUCHPLBPRIO  =>  TIEC440ICURDTOUCHPLBPRIO_indelay,
	TIEC440PIR  =>  TIEC440PIR_indelay,
	TIEC440PVR  =>  TIEC440PVR_indelay,
	TIEC440USERRESET  =>  TIEC440USERRESET_indelay,
	TIEDCRBASEADDR  =>  TIEDCRBASEADDR_indelay,
	TRCC440TRACEDISABLE  =>  TRCC440TRACEDISABLE_indelay,
	TRCC440TRIGGEREVENTIN  =>  TRCC440TRIGGEREVENTIN_indelay
	);

	INIPROC : process
	begin
       case PPCS0_WIDTH_128N64 is
           when FALSE   =>  PPCS0_WIDTH_128N64_BINARY <= '0';
           when TRUE    =>  PPCS0_WIDTH_128N64_BINARY <= '1';
           when others  =>  assert FALSE report "Error : PPCS0_WIDTH_128N64 is neither TRUE nor FALSE." severity error;
       end case;
       case PPCS1_WIDTH_128N64 is
           when FALSE   =>  PPCS1_WIDTH_128N64_BINARY <= '0';
           when TRUE    =>  PPCS1_WIDTH_128N64_BINARY <= '1';
           when others  =>  assert FALSE report "Error : PPCS1_WIDTH_128N64 is neither TRUE nor FALSE." severity error;
       end case;
       case PPCDM_ASYNCMODE is
           when FALSE   =>  PPCDM_ASYNCMODE_BINARY <= '0';
           when TRUE    =>  PPCDM_ASYNCMODE_BINARY <= '1';
           when others  =>  assert FALSE report "Error : PPCDM_ASYNCMODE is neither TRUE nor FALSE." severity error;
       end case;
       case PPCDS_ASYNCMODE is
           when FALSE   =>  PPCDS_ASYNCMODE_BINARY <= '0';
           when TRUE    =>  PPCDS_ASYNCMODE_BINARY <= '1';
           when others  =>  assert FALSE report "Error : PPCDS_ASYNCMODE is neither TRUE nor FALSE." severity error;
       end case;
       case DCR_AUTOLOCK_ENABLE is
           when FALSE   =>  DCR_AUTOLOCK_ENABLE_BINARY <= '0';
           when TRUE    =>  DCR_AUTOLOCK_ENABLE_BINARY <= '1';
           when others  =>  assert FALSE report "Error : DCR_AUTOLOCK_ENABLE is neither TRUE nor FALSE." severity error;
       end case;
       case CLOCK_DELAY is
--           when FALSE   =>  CLOCK_DELAY_BINARY <= "00100";
           when FALSE   =>  CLOCK_DELAY_BINARY <= "10000";
           when TRUE    =>  CLOCK_DELAY_BINARY <= "00000";
           when others  =>  assert FALSE report "Error : CLOCK_DELAY is neither TRUE nor FALSE." severity error;
       end case;
	wait;
	end process INIPROC;

	TIMING : process

	variable Tmkr_CPMC440CORECLOCKINACTIVE_JTGC440TCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_CPMINTERCONNECTCLKNTO1_CPMINTERCONNECTCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DBGC440DEBUGHALT_CPMC440CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DBGC440SYSTEMSTATUS0_JTGC440TCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DBGC440SYSTEMSTATUS1_JTGC440TCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DBGC440SYSTEMSTATUS2_JTGC440TCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DBGC440SYSTEMSTATUS3_JTGC440TCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DBGC440SYSTEMSTATUS4_JTGC440TCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DBGC440UNCONDDEBUGEVENT_CPMC440CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMACK_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN0_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN10_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN11_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN12_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN13_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN14_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN15_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN16_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN17_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN18_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN19_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN1_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN20_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN21_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN22_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN23_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN24_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN25_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN26_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN27_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN28_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN29_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN2_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN30_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN31_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN3_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN4_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN5_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN6_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN7_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN8_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMDBUSIN9_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDMTIMEOUTWAIT_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSABUS0_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSABUS1_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSABUS2_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSABUS3_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSABUS4_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSABUS5_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSABUS6_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSABUS7_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSABUS8_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSABUS9_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT0_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT10_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT11_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT12_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT13_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT14_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT15_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT16_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT17_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT18_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT19_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT1_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT20_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT21_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT22_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT23_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT24_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT25_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT26_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT27_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT28_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT29_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT2_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT30_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT31_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT3_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT4_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT5_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT6_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT7_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT8_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSDBUSOUT9_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSREAD_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_DCRPPCDSWRITE_CPMDCRCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUCONFIRMINSTR_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUCR0_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUCR1_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUCR2_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUCR3_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUDONE_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUEXCEPTION_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUFPSCRFEX_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT0_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT10_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT11_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT12_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT13_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT14_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT15_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT16_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT17_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT18_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT19_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT1_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT20_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT21_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT22_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT23_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT24_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT25_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT26_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT27_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT28_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT29_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT2_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT30_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT31_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT3_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT4_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT5_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT6_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT7_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT8_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULT9_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPURESULTVALID_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSLEEPNOTREADY_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA0_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA100_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA101_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA102_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA103_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA104_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA105_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA106_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA107_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA108_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA109_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA10_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA110_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA111_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA112_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA113_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA114_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA115_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA116_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA117_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA118_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA119_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA11_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA120_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA121_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA122_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA123_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA124_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA125_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA126_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA127_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA12_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA13_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA14_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA15_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA16_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA17_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA18_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA19_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA1_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA20_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA21_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA22_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA23_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA24_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA25_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA26_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA27_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA28_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA29_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA2_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA30_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA31_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA32_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA33_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA34_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA35_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA36_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA37_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA38_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA39_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA3_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA40_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA41_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA42_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA43_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA44_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA45_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA46_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA47_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA48_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA49_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA4_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA50_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA51_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA52_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA53_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA54_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA55_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA56_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA57_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA58_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA59_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA5_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA60_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA61_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA62_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA63_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA64_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA65_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA66_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA67_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA68_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA69_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA6_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA70_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA71_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA72_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA73_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA74_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA75_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA76_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA77_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA78_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA79_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA7_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA80_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA81_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA82_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA83_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA84_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA85_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA86_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA87_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA88_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA89_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA8_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA90_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA91_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA92_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA93_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA94_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA95_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA96_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA97_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA98_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA99_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_FCMAPUSTOREDATA9_CPMFCMCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_JTGC440TDI_JTGC440TCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_JTGC440TMS_JTGC440TCK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RSTENGINEREQ_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD0_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD10_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD11_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD12_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD13_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD14_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD15_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD16_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD17_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD18_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD19_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD1_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD20_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD21_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD22_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD23_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD24_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD25_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD26_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD27_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD28_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD29_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD2_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD30_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD31_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD3_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD4_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD5_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD6_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD7_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD8_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXD9_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXEOFN_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXEOPN_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXREM0_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXREM1_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXREM2_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXREM3_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXSOFN_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXSOPN_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0RXSRCRDYN_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA0TXDSTRDYN_CPMDMA0LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RSTENGINEREQ_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD0_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD10_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD11_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD12_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD13_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD14_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD15_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD16_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD17_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD18_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD19_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD1_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD20_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD21_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD22_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD23_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD24_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD25_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD26_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD27_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD28_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD29_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD2_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD30_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD31_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD3_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD4_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD5_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD6_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD7_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD8_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXD9_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXEOFN_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXEOPN_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXREM0_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXREM1_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXREM2_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXREM3_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXSOFN_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXSOPN_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1RXSRCRDYN_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA1TXDSTRDYN_CPMDMA1LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RSTENGINEREQ_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD0_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD10_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD11_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD12_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD13_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD14_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD15_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD16_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD17_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD18_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD19_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD1_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD20_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD21_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD22_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD23_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD24_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD25_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD26_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD27_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD28_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD29_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD2_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD30_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD31_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD3_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD4_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD5_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD6_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD7_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD8_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXD9_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXEOFN_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXEOPN_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXREM0_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXREM1_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXREM2_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXREM3_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXSOFN_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXSOPN_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2RXSRCRDYN_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA2TXDSTRDYN_CPMDMA2LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RSTENGINEREQ_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD0_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD10_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD11_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD12_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD13_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD14_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD15_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD16_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD17_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD18_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD19_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD1_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD20_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD21_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD22_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD23_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD24_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD25_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD26_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD27_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD28_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD29_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD2_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD30_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD31_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD3_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD4_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD5_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD6_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD7_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD8_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXD9_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXEOFN_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXEOPN_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXREM0_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXREM1_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXREM2_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXREM3_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXSOFN_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXSOPN_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3RXSRCRDYN_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_LLDMA3TXDSTRDYN_CPMDMA3LLCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIADDRREADYTOACCEPT_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA0_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA100_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA101_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA102_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA103_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA104_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA105_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA106_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA107_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA108_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA109_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA10_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA110_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA111_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA112_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA113_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA114_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA115_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA116_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA117_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA118_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA119_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA11_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA120_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA121_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA122_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA123_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA124_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA125_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA126_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA127_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA12_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA13_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA14_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA15_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA16_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA17_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA18_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA19_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA1_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA20_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA21_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA22_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA23_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA24_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA25_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA26_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA27_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA28_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA29_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA2_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA30_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA31_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA32_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA33_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA34_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA35_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA36_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA37_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA38_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA39_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA3_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA40_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA41_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA42_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA43_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA44_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA45_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA46_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA47_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA48_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA49_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA4_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA50_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA51_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA52_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA53_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA54_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA55_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA56_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA57_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA58_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA59_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA5_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA60_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA61_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA62_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA63_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA64_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA65_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA66_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA67_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA68_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA69_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA6_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA70_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA71_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA72_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA73_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA74_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA75_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA76_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA77_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA78_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA79_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA7_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA80_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA81_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA82_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA83_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA84_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA85_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA86_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA87_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA88_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA89_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA8_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA90_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA91_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA92_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA93_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA94_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA95_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA96_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA97_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA98_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA99_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATA9_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATAERR_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_MCMIREADDATAVALID_CPMMCCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMADDRACK_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMMBUSY_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMMIRQ_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMMRDERR_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMMWRERR_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDBTERM_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDACK_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS0_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS100_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS101_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS102_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS103_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS104_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS105_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS106_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS107_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS108_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS109_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS10_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS110_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS111_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS112_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS113_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS114_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS115_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS116_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS117_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS118_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS119_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS11_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS120_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS121_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS122_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS123_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS124_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS125_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS126_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS127_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS12_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS13_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS14_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS15_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS16_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS17_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS18_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS19_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS1_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS20_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS21_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS22_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS23_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS24_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS25_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS26_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS27_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS28_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS29_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS2_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS30_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS31_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS32_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS33_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS34_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS35_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS36_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS37_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS38_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS39_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS3_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS40_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS41_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS42_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS43_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS44_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS45_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS46_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS47_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS48_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS49_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS4_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS50_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS51_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS52_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS53_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS54_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS55_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS56_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS57_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS58_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS59_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS5_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS60_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS61_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS62_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS63_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS64_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS65_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS66_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS67_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS68_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS69_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS6_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS70_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS71_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS72_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS73_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS74_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS75_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS76_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS77_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS78_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS79_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS7_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS80_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS81_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS82_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS83_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS84_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS85_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS86_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS87_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS88_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS89_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS8_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS90_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS91_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS92_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS93_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS94_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS95_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS96_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS97_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS98_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS99_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDDBUS9_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDPENDPRI0_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDPENDPRI1_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDPENDREQ_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDWDADDR0_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDWDADDR1_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDWDADDR2_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMRDWDADDR3_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMREARBITRATE_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMREQPRI0_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMREQPRI1_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMSSIZE0_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMSSIZE1_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMTIMEOUT_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMWRBTERM_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMWRDACK_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMWRPENDPRI0_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMWRPENDPRI1_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCMWRPENDREQ_CPMPPCMPLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABORT_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS0_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS10_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS11_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS12_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS13_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS14_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS15_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS16_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS17_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS18_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS19_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS1_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS20_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS21_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS22_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS23_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS24_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS25_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS26_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS27_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS28_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS29_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS2_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS30_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS31_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS3_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS4_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS5_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS6_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS7_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS8_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0ABUS9_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE0_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE10_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE11_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE12_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE13_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE14_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE15_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE1_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE2_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE3_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE4_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE5_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE6_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE7_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE8_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BE9_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0BUSLOCK_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0LOCKERR_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0MASTERID0_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0MASTERID1_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0MSIZE0_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0MSIZE1_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0PAVALID_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0RDBURST_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0RDPENDPRI0_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0RDPENDPRI1_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0RDPENDREQ_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0RDPRIM_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0REQPRI0_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0REQPRI1_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0RNW_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0SAVALID_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0SIZE0_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0SIZE1_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0SIZE2_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0SIZE3_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE0_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE10_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE11_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE12_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE13_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE14_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE15_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE1_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE2_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE3_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE4_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE5_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE6_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE7_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE8_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TATTRIBUTE9_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TYPE0_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TYPE1_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0TYPE2_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0UABUS28_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0UABUS29_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0UABUS30_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0UABUS31_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRBURST_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS0_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS100_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS101_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS102_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS103_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS104_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS105_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS106_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS107_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS108_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS109_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS10_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS110_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS111_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS112_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS113_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS114_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS115_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS116_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS117_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS118_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS119_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS11_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS120_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS121_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS122_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS123_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS124_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS125_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS126_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS127_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS12_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS13_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS14_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS15_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS16_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS17_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS18_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS19_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS1_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS20_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS21_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS22_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS23_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS24_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS25_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS26_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS27_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS28_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS29_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS2_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS30_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS31_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS32_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS33_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS34_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS35_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS36_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS37_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS38_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS39_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS3_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS40_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS41_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS42_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS43_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS44_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS45_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS46_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS47_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS48_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS49_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS4_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS50_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS51_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS52_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS53_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS54_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS55_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS56_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS57_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS58_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS59_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS5_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS60_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS61_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS62_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS63_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS64_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS65_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS66_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS67_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS68_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS69_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS6_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS70_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS71_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS72_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS73_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS74_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS75_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS76_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS77_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS78_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS79_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS7_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS80_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS81_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS82_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS83_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS84_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS85_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS86_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS87_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS88_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS89_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS8_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS90_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS91_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS92_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS93_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS94_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS95_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS96_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS97_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS98_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS99_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRDBUS9_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRPENDPRI0_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRPENDPRI1_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRPENDREQ_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS0WRPRIM_CPMPPCS0PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABORT_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS0_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS10_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS11_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS12_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS13_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS14_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS15_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS16_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS17_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS18_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS19_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS1_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS20_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS21_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS22_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS23_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS24_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS25_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS26_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS27_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS28_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS29_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS2_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS30_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS31_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS3_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS4_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS5_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS6_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS7_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS8_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1ABUS9_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE0_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE10_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE11_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE12_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE13_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE14_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE15_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE1_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE2_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE3_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE4_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE5_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE6_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE7_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE8_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BE9_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1BUSLOCK_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1LOCKERR_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1MASTERID0_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1MASTERID1_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1MSIZE0_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1MSIZE1_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1PAVALID_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1RDBURST_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1RDPENDPRI0_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1RDPENDPRI1_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1RDPENDREQ_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1RDPRIM_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1REQPRI0_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1REQPRI1_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1RNW_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1SAVALID_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1SIZE0_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1SIZE1_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1SIZE2_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1SIZE3_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE0_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE10_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE11_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE12_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE13_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE14_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE15_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE1_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE2_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE3_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE4_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE5_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE6_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE7_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE8_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TATTRIBUTE9_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TYPE0_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TYPE1_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1TYPE2_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1UABUS28_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1UABUS29_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1UABUS30_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1UABUS31_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRBURST_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS0_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS100_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS101_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS102_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS103_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS104_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS105_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS106_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS107_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS108_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS109_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS10_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS110_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS111_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS112_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS113_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS114_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS115_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS116_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS117_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS118_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS119_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS11_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS120_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS121_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS122_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS123_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS124_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS125_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS126_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS127_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS12_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS13_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS14_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS15_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS16_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS17_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS18_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS19_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS1_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS20_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS21_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS22_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS23_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS24_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS25_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS26_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS27_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS28_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS29_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS2_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS30_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS31_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS32_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS33_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS34_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS35_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS36_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS37_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS38_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS39_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS3_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS40_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS41_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS42_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS43_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS44_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS45_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS46_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS47_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS48_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS49_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS4_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS50_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS51_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS52_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS53_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS54_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS55_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS56_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS57_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS58_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS59_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS5_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS60_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS61_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS62_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS63_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS64_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS65_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS66_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS67_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS68_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS69_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS6_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS70_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS71_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS72_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS73_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS74_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS75_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS76_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS77_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS78_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS79_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS7_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS80_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS81_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS82_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS83_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS84_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS85_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS86_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS87_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS88_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS89_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS8_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS90_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS91_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS92_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS93_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS94_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS95_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS96_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS97_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS98_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS99_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRDBUS9_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRPENDPRI0_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRPENDPRI1_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRPENDREQ_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_PLBPPCS1WRPRIM_CPMPPCS1PLBCLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_TRCC440TRACEDISABLE_CPMC440CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tmkr_TRCC440TRIGGEREVENTIN_CPMC440CLK_posedge : VitalTimingDataType := VitalTimingDataInit;
	variable Tviol_CPMC440CORECLOCKINACTIVE_JTGC440TCK_posedge : STD_ULOGIC := '0';
	variable Tviol_CPMINTERCONNECTCLKNTO1_CPMINTERCONNECTCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DBGC440DEBUGHALT_CPMC440CLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DBGC440SYSTEMSTATUS0_JTGC440TCK_posedge : STD_ULOGIC := '0';
	variable Tviol_DBGC440SYSTEMSTATUS1_JTGC440TCK_posedge : STD_ULOGIC := '0';
	variable Tviol_DBGC440SYSTEMSTATUS2_JTGC440TCK_posedge : STD_ULOGIC := '0';
	variable Tviol_DBGC440SYSTEMSTATUS3_JTGC440TCK_posedge : STD_ULOGIC := '0';
	variable Tviol_DBGC440SYSTEMSTATUS4_JTGC440TCK_posedge : STD_ULOGIC := '0';
	variable Tviol_DBGC440UNCONDDEBUGEVENT_CPMC440CLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMACK_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN0_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN10_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN11_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN12_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN13_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN14_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN15_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN16_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN17_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN18_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN19_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN1_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN20_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN21_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN22_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN23_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN24_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN25_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN26_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN27_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN28_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN29_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN2_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN30_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN31_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN3_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN4_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN5_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN6_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN7_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN8_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMDBUSIN9_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDMTIMEOUTWAIT_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSABUS0_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSABUS1_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSABUS2_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSABUS3_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSABUS4_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSABUS5_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSABUS6_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSABUS7_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSABUS8_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSABUS9_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT0_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT10_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT11_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT12_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT13_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT14_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT15_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT16_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT17_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT18_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT19_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT1_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT20_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT21_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT22_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT23_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT24_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT25_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT26_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT27_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT28_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT29_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT2_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT30_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT31_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT3_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT4_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT5_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT6_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT7_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT8_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSDBUSOUT9_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSREAD_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_DCRPPCDSWRITE_CPMDCRCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUCONFIRMINSTR_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUCR0_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUCR1_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUCR2_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUCR3_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUDONE_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUEXCEPTION_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUFPSCRFEX_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT0_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT10_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT11_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT12_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT13_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT14_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT15_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT16_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT17_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT18_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT19_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT1_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT20_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT21_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT22_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT23_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT24_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT25_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT26_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT27_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT28_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT29_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT2_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT30_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT31_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT3_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT4_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT5_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT6_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT7_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT8_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULT9_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPURESULTVALID_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSLEEPNOTREADY_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA0_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA100_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA101_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA102_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA103_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA104_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA105_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA106_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA107_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA108_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA109_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA10_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA110_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA111_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA112_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA113_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA114_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA115_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA116_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA117_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA118_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA119_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA11_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA120_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA121_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA122_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA123_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA124_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA125_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA126_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA127_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA12_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA13_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA14_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA15_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA16_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA17_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA18_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA19_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA1_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA20_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA21_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA22_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA23_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA24_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA25_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA26_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA27_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA28_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA29_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA2_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA30_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA31_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA32_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA33_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA34_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA35_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA36_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA37_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA38_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA39_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA3_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA40_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA41_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA42_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA43_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA44_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA45_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA46_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA47_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA48_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA49_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA4_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA50_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA51_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA52_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA53_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA54_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA55_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA56_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA57_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA58_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA59_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA5_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA60_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA61_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA62_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA63_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA64_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA65_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA66_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA67_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA68_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA69_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA6_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA70_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA71_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA72_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA73_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA74_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA75_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA76_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA77_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA78_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA79_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA7_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA80_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA81_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA82_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA83_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA84_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA85_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA86_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA87_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA88_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA89_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA8_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA90_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA91_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA92_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA93_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA94_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA95_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA96_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA97_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA98_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA99_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_FCMAPUSTOREDATA9_CPMFCMCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_JTGC440TDI_JTGC440TCK_posedge : STD_ULOGIC := '0';
	variable Tviol_JTGC440TMS_JTGC440TCK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RSTENGINEREQ_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD0_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD10_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD11_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD12_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD13_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD14_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD15_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD16_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD17_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD18_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD19_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD1_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD20_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD21_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD22_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD23_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD24_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD25_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD26_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD27_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD28_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD29_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD2_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD30_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD31_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD3_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD4_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD5_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD6_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD7_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD8_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXD9_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXEOFN_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXEOPN_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXREM0_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXREM1_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXREM2_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXREM3_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXSOFN_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXSOPN_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0RXSRCRDYN_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA0TXDSTRDYN_CPMDMA0LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RSTENGINEREQ_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD0_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD10_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD11_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD12_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD13_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD14_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD15_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD16_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD17_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD18_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD19_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD1_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD20_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD21_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD22_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD23_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD24_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD25_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD26_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD27_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD28_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD29_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD2_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD30_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD31_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD3_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD4_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD5_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD6_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD7_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD8_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXD9_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXEOFN_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXEOPN_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXREM0_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXREM1_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXREM2_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXREM3_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXSOFN_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXSOPN_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1RXSRCRDYN_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA1TXDSTRDYN_CPMDMA1LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RSTENGINEREQ_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD0_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD10_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD11_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD12_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD13_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD14_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD15_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD16_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD17_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD18_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD19_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD1_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD20_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD21_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD22_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD23_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD24_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD25_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD26_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD27_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD28_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD29_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD2_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD30_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD31_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD3_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD4_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD5_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD6_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD7_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD8_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXD9_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXEOFN_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXEOPN_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXREM0_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXREM1_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXREM2_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXREM3_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXSOFN_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXSOPN_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2RXSRCRDYN_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA2TXDSTRDYN_CPMDMA2LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RSTENGINEREQ_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD0_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD10_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD11_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD12_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD13_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD14_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD15_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD16_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD17_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD18_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD19_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD1_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD20_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD21_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD22_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD23_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD24_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD25_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD26_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD27_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD28_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD29_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD2_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD30_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD31_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD3_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD4_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD5_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD6_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD7_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD8_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXD9_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXEOFN_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXEOPN_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXREM0_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXREM1_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXREM2_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXREM3_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXSOFN_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXSOPN_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3RXSRCRDYN_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_LLDMA3TXDSTRDYN_CPMDMA3LLCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIADDRREADYTOACCEPT_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA0_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA100_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA101_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA102_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA103_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA104_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA105_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA106_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA107_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA108_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA109_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA10_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA110_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA111_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA112_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA113_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA114_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA115_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA116_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA117_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA118_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA119_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA11_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA120_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA121_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA122_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA123_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA124_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA125_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA126_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA127_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA12_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA13_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA14_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA15_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA16_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA17_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA18_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA19_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA1_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA20_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA21_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA22_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA23_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA24_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA25_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA26_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA27_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA28_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA29_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA2_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA30_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA31_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA32_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA33_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA34_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA35_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA36_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA37_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA38_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA39_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA3_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA40_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA41_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA42_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA43_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA44_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA45_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA46_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA47_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA48_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA49_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA4_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA50_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA51_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA52_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA53_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA54_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA55_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA56_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA57_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA58_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA59_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA5_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA60_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA61_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA62_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA63_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA64_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA65_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA66_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA67_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA68_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA69_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA6_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA70_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA71_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA72_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA73_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA74_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA75_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA76_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA77_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA78_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA79_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA7_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA80_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA81_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA82_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA83_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA84_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA85_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA86_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA87_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA88_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA89_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA8_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA90_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA91_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA92_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA93_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA94_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA95_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA96_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA97_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA98_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA99_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATA9_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATAERR_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_MCMIREADDATAVALID_CPMMCCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMADDRACK_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMMBUSY_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMMIRQ_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMMRDERR_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMMWRERR_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDBTERM_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDACK_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS0_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS100_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS101_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS102_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS103_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS104_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS105_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS106_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS107_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS108_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS109_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS10_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS110_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS111_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS112_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS113_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS114_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS115_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS116_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS117_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS118_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS119_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS11_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS120_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS121_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS122_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS123_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS124_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS125_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS126_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS127_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS12_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS13_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS14_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS15_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS16_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS17_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS18_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS19_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS1_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS20_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS21_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS22_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS23_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS24_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS25_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS26_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS27_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS28_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS29_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS2_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS30_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS31_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS32_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS33_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS34_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS35_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS36_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS37_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS38_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS39_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS3_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS40_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS41_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS42_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS43_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS44_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS45_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS46_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS47_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS48_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS49_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS4_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS50_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS51_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS52_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS53_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS54_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS55_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS56_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS57_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS58_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS59_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS5_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS60_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS61_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS62_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS63_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS64_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS65_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS66_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS67_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS68_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS69_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS6_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS70_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS71_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS72_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS73_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS74_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS75_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS76_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS77_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS78_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS79_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS7_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS80_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS81_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS82_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS83_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS84_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS85_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS86_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS87_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS88_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS89_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS8_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS90_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS91_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS92_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS93_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS94_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS95_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS96_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS97_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS98_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS99_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDDBUS9_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDPENDPRI0_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDPENDPRI1_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDPENDREQ_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDWDADDR0_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDWDADDR1_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDWDADDR2_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMRDWDADDR3_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMREARBITRATE_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMREQPRI0_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMREQPRI1_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMSSIZE0_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMSSIZE1_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMTIMEOUT_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMWRBTERM_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMWRDACK_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMWRPENDPRI0_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMWRPENDPRI1_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCMWRPENDREQ_CPMPPCMPLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABORT_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS0_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS10_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS11_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS12_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS13_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS14_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS15_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS16_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS17_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS18_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS19_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS1_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS20_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS21_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS22_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS23_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS24_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS25_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS26_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS27_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS28_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS29_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS2_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS30_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS31_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS3_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS4_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS5_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS6_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS7_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS8_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0ABUS9_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE0_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE10_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE11_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE12_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE13_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE14_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE15_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE1_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE2_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE3_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE4_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE5_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE6_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE7_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE8_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BE9_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0BUSLOCK_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0LOCKERR_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0MASTERID0_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0MASTERID1_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0MSIZE0_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0MSIZE1_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0PAVALID_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0RDBURST_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0RDPENDPRI0_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0RDPENDPRI1_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0RDPENDREQ_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0RDPRIM_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0REQPRI0_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0REQPRI1_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0RNW_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0SAVALID_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0SIZE0_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0SIZE1_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0SIZE2_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0SIZE3_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE0_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE10_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE11_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE12_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE13_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE14_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE15_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE1_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE2_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE3_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE4_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE5_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE6_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE7_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE8_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TATTRIBUTE9_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TYPE0_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TYPE1_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0TYPE2_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0UABUS28_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0UABUS29_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0UABUS30_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0UABUS31_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRBURST_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS0_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS100_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS101_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS102_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS103_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS104_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS105_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS106_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS107_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS108_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS109_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS10_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS110_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS111_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS112_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS113_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS114_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS115_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS116_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS117_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS118_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS119_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS11_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS120_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS121_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS122_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS123_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS124_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS125_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS126_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS127_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS12_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS13_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS14_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS15_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS16_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS17_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS18_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS19_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS1_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS20_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS21_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS22_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS23_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS24_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS25_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS26_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS27_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS28_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS29_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS2_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS30_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS31_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS32_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS33_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS34_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS35_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS36_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS37_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS38_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS39_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS3_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS40_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS41_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS42_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS43_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS44_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS45_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS46_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS47_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS48_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS49_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS4_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS50_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS51_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS52_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS53_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS54_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS55_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS56_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS57_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS58_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS59_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS5_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS60_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS61_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS62_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS63_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS64_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS65_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS66_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS67_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS68_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS69_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS6_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS70_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS71_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS72_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS73_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS74_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS75_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS76_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS77_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS78_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS79_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS7_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS80_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS81_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS82_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS83_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS84_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS85_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS86_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS87_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS88_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS89_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS8_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS90_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS91_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS92_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS93_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS94_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS95_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS96_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS97_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS98_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS99_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRDBUS9_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRPENDPRI0_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRPENDPRI1_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRPENDREQ_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS0WRPRIM_CPMPPCS0PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABORT_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS0_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS10_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS11_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS12_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS13_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS14_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS15_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS16_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS17_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS18_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS19_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS1_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS20_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS21_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS22_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS23_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS24_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS25_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS26_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS27_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS28_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS29_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS2_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS30_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS31_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS3_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS4_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS5_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS6_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS7_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS8_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1ABUS9_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE0_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE10_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE11_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE12_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE13_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE14_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE15_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE1_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE2_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE3_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE4_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE5_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE6_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE7_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE8_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BE9_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1BUSLOCK_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1LOCKERR_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1MASTERID0_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1MASTERID1_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1MSIZE0_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1MSIZE1_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1PAVALID_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1RDBURST_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1RDPENDPRI0_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1RDPENDPRI1_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1RDPENDREQ_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1RDPRIM_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1REQPRI0_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1REQPRI1_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1RNW_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1SAVALID_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1SIZE0_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1SIZE1_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1SIZE2_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1SIZE3_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE0_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE10_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE11_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE12_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE13_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE14_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE15_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE1_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE2_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE3_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE4_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE5_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE6_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE7_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE8_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TATTRIBUTE9_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TYPE0_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TYPE1_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1TYPE2_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1UABUS28_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1UABUS29_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1UABUS30_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1UABUS31_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRBURST_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS0_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS100_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS101_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS102_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS103_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS104_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS105_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS106_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS107_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS108_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS109_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS10_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS110_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS111_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS112_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS113_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS114_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS115_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS116_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS117_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS118_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS119_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS11_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS120_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS121_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS122_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS123_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS124_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS125_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS126_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS127_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS12_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS13_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS14_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS15_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS16_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS17_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS18_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS19_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS1_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS20_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS21_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS22_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS23_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS24_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS25_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS26_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS27_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS28_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS29_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS2_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS30_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS31_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS32_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS33_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS34_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS35_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS36_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS37_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS38_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS39_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS3_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS40_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS41_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS42_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS43_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS44_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS45_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS46_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS47_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS48_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS49_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS4_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS50_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS51_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS52_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS53_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS54_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS55_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS56_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS57_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS58_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS59_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS5_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS60_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS61_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS62_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS63_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS64_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS65_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS66_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS67_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS68_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS69_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS6_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS70_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS71_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS72_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS73_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS74_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS75_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS76_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS77_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS78_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS79_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS7_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS80_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS81_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS82_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS83_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS84_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS85_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS86_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS87_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS88_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS89_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS8_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS90_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS91_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS92_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS93_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS94_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS95_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS96_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS97_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS98_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS99_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRDBUS9_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRPENDPRI0_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRPENDPRI1_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRPENDREQ_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_PLBPPCS1WRPRIM_CPMPPCS1PLBCLK_posedge : STD_ULOGIC := '0';
	variable Tviol_TRCC440TRACEDISABLE_CPMC440CLK_posedge : STD_ULOGIC := '0';
	variable Tviol_TRCC440TRIGGEREVENTIN_CPMC440CLK_posedge : STD_ULOGIC := '0';

	variable  DMA0LLRSTENGINEACK_GlitchData : VitalGlitchDataType;
	variable  DMA0LLRXDSTRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD0_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD1_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD2_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD3_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD4_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD5_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD6_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD7_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD8_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD9_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD10_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD11_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD12_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD13_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD14_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD15_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD16_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD17_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD18_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD19_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD20_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD21_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD22_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD23_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD24_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD25_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD26_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD27_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD28_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD29_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD30_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXD31_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXEOFN_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXEOPN_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXREM0_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXREM1_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXREM2_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXREM3_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXSOFN_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXSOPN_GlitchData : VitalGlitchDataType;
	variable  DMA0LLTXSRCRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA0RXIRQ_GlitchData : VitalGlitchDataType;
	variable  DMA0TXIRQ_GlitchData : VitalGlitchDataType;
	variable  DMA1LLRSTENGINEACK_GlitchData : VitalGlitchDataType;
	variable  DMA1LLRXDSTRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD0_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD1_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD2_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD3_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD4_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD5_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD6_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD7_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD8_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD9_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD10_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD11_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD12_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD13_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD14_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD15_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD16_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD17_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD18_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD19_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD20_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD21_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD22_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD23_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD24_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD25_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD26_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD27_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD28_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD29_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD30_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXD31_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXEOFN_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXEOPN_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXREM0_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXREM1_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXREM2_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXREM3_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXSOFN_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXSOPN_GlitchData : VitalGlitchDataType;
	variable  DMA1LLTXSRCRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA1RXIRQ_GlitchData : VitalGlitchDataType;
	variable  DMA1TXIRQ_GlitchData : VitalGlitchDataType;
	variable  DMA2LLRSTENGINEACK_GlitchData : VitalGlitchDataType;
	variable  DMA2LLRXDSTRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD0_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD1_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD2_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD3_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD4_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD5_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD6_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD7_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD8_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD9_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD10_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD11_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD12_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD13_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD14_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD15_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD16_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD17_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD18_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD19_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD20_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD21_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD22_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD23_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD24_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD25_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD26_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD27_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD28_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD29_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD30_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXD31_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXEOFN_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXEOPN_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXREM0_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXREM1_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXREM2_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXREM3_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXSOFN_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXSOPN_GlitchData : VitalGlitchDataType;
	variable  DMA2LLTXSRCRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA2RXIRQ_GlitchData : VitalGlitchDataType;
	variable  DMA2TXIRQ_GlitchData : VitalGlitchDataType;
	variable  DMA3LLRSTENGINEACK_GlitchData : VitalGlitchDataType;
	variable  DMA3LLRXDSTRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD0_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD1_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD2_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD3_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD4_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD5_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD6_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD7_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD8_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD9_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD10_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD11_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD12_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD13_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD14_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD15_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD16_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD17_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD18_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD19_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD20_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD21_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD22_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD23_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD24_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD25_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD26_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD27_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD28_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD29_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD30_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXD31_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXEOFN_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXEOPN_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXREM0_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXREM1_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXREM2_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXREM3_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXSOFN_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXSOPN_GlitchData : VitalGlitchDataType;
	variable  DMA3LLTXSRCRDYN_GlitchData : VitalGlitchDataType;
	variable  DMA3RXIRQ_GlitchData : VitalGlitchDataType;
	variable  DMA3TXIRQ_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS0_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS1_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS2_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS3_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS4_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS5_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS6_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS7_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS8_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRABUS9_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT0_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT1_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT2_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT3_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT4_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT5_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT6_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT7_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT8_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT9_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT10_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT11_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT12_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT13_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT14_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT15_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT16_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT17_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT18_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT19_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT20_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT21_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT22_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT23_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT24_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT25_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT26_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT27_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT28_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT29_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT30_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRDBUSOUT31_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRREAD_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRUABUS20_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRUABUS21_GlitchData : VitalGlitchDataType;
	variable  PPCDMDCRWRITE_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABORT_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS0_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS1_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS2_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS3_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS4_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS5_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS6_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS7_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS8_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS9_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS10_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS11_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS12_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS13_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS14_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS15_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS16_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS17_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS18_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS19_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS20_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS21_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS22_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS23_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS24_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS25_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS26_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS27_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS28_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS29_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS30_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBABUS31_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE0_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE1_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE2_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE3_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE4_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE5_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE6_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE7_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE8_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE9_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE10_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE11_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE12_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE13_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE14_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBE15_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBBUSLOCK_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBLOCKERR_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBPRIORITY0_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBPRIORITY1_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBRDBURST_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBREQUEST_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBRNW_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBSIZE0_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBSIZE1_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBSIZE2_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBSIZE3_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE0_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE1_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE2_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE3_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE4_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE5_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE6_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE7_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE8_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE9_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE10_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE11_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE12_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE13_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE14_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTATTRIBUTE15_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTYPE0_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTYPE1_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBTYPE2_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBUABUS28_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBUABUS29_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBUABUS30_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBUABUS31_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRBURST_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS0_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS1_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS2_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS3_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS4_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS5_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS6_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS7_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS8_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS9_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS10_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS11_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS12_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS13_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS14_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS15_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS16_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS17_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS18_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS19_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS20_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS21_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS22_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS23_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS24_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS25_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS26_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS27_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS28_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS29_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS30_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS31_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS32_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS33_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS34_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS35_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS36_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS37_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS38_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS39_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS40_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS41_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS42_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS43_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS44_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS45_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS46_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS47_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS48_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS49_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS50_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS51_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS52_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS53_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS54_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS55_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS56_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS57_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS58_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS59_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS60_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS61_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS62_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS63_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS64_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS65_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS66_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS67_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS68_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS69_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS70_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS71_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS72_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS73_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS74_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS75_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS76_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS77_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS78_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS79_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS80_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS81_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS82_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS83_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS84_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS85_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS86_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS87_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS88_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS89_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS90_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS91_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS92_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS93_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS94_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS95_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS96_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS97_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS98_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS99_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS100_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS101_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS102_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS103_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS104_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS105_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS106_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS107_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS108_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS109_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS110_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS111_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS112_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS113_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS114_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS115_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS116_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS117_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS118_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS119_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS120_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS121_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS122_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS123_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS124_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS125_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS126_GlitchData : VitalGlitchDataType;
	variable  PPCMPLBWRDBUS127_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBADDRACK_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMBUSY0_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMBUSY1_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMBUSY2_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMBUSY3_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMIRQ0_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMIRQ1_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMIRQ2_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMIRQ3_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMRDERR0_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMRDERR1_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMRDERR2_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMRDERR3_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMWRERR0_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMWRERR1_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMWRERR2_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBMWRERR3_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDBTERM_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDCOMP_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDACK_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS0_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS1_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS2_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS3_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS4_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS5_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS6_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS7_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS8_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS9_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS10_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS11_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS12_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS13_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS14_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS15_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS16_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS17_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS18_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS19_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS20_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS21_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS22_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS23_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS24_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS25_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS26_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS27_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS28_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS29_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS30_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS31_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS32_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS33_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS34_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS35_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS36_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS37_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS38_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS39_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS40_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS41_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS42_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS43_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS44_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS45_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS46_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS47_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS48_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS49_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS50_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS51_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS52_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS53_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS54_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS55_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS56_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS57_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS58_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS59_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS60_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS61_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS62_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS63_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS64_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS65_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS66_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS67_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS68_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS69_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS70_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS71_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS72_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS73_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS74_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS75_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS76_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS77_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS78_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS79_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS80_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS81_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS82_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS83_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS84_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS85_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS86_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS87_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS88_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS89_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS90_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS91_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS92_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS93_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS94_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS95_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS96_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS97_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS98_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS99_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS100_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS101_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS102_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS103_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS104_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS105_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS106_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS107_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS108_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS109_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS110_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS111_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS112_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS113_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS114_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS115_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS116_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS117_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS118_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS119_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS120_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS121_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS122_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS123_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS124_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS125_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS126_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDDBUS127_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDWDADDR0_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDWDADDR1_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDWDADDR2_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBRDWDADDR3_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBREARBITRATE_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBSSIZE0_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBSSIZE1_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBWAIT_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBWRBTERM_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBWRCOMP_GlitchData : VitalGlitchDataType;
	variable  PPCS0PLBWRDACK_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBADDRACK_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMBUSY0_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMBUSY1_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMBUSY2_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMBUSY3_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMIRQ0_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMIRQ1_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMIRQ2_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMIRQ3_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMRDERR0_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMRDERR1_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMRDERR2_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMRDERR3_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMWRERR0_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMWRERR1_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMWRERR2_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBMWRERR3_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDBTERM_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDCOMP_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDACK_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS0_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS1_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS2_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS3_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS4_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS5_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS6_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS7_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS8_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS9_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS10_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS11_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS12_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS13_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS14_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS15_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS16_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS17_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS18_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS19_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS20_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS21_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS22_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS23_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS24_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS25_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS26_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS27_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS28_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS29_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS30_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS31_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS32_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS33_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS34_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS35_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS36_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS37_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS38_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS39_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS40_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS41_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS42_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS43_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS44_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS45_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS46_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS47_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS48_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS49_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS50_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS51_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS52_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS53_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS54_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS55_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS56_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS57_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS58_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS59_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS60_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS61_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS62_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS63_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS64_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS65_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS66_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS67_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS68_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS69_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS70_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS71_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS72_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS73_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS74_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS75_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS76_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS77_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS78_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS79_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS80_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS81_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS82_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS83_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS84_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS85_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS86_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS87_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS88_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS89_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS90_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS91_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS92_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS93_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS94_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS95_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS96_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS97_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS98_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS99_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS100_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS101_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS102_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS103_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS104_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS105_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS106_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS107_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS108_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS109_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS110_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS111_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS112_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS113_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS114_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS115_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS116_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS117_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS118_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS119_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS120_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS121_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS122_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS123_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS124_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS125_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS126_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDDBUS127_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDWDADDR0_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDWDADDR1_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDWDADDR2_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBRDWDADDR3_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBREARBITRATE_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBSSIZE0_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBSSIZE1_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBWAIT_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBWRBTERM_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBWRCOMP_GlitchData : VitalGlitchDataType;
	variable  PPCS1PLBWRDACK_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECFPUOP_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECLDSTXFERSIZE0_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECLDSTXFERSIZE1_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECLDSTXFERSIZE2_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECLOAD_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECNONAUTON_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECSTORE_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECUDI0_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECUDI1_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECUDI2_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECUDI3_GlitchData : VitalGlitchDataType;
	variable  APUFCMDECUDIVALID_GlitchData : VitalGlitchDataType;
	variable  APUFCMENDIAN_GlitchData : VitalGlitchDataType;
	variable  APUFCMFLUSH_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION0_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION1_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION2_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION3_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION4_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION5_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION6_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION7_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION8_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION9_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION10_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION11_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION12_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION13_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION14_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION15_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION16_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION17_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION18_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION19_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION20_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION21_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION22_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION23_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION24_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION25_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION26_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION27_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION28_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION29_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION30_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRUCTION31_GlitchData : VitalGlitchDataType;
	variable  APUFCMINSTRVALID_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADBYTEADDR0_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADBYTEADDR1_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADBYTEADDR2_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADBYTEADDR3_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA0_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA1_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA2_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA3_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA4_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA5_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA6_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA7_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA8_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA9_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA10_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA11_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA12_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA13_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA14_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA15_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA16_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA17_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA18_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA19_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA20_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA21_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA22_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA23_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA24_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA25_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA26_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA27_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA28_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA29_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA30_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA31_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA32_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA33_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA34_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA35_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA36_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA37_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA38_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA39_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA40_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA41_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA42_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA43_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA44_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA45_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA46_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA47_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA48_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA49_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA50_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA51_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA52_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA53_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA54_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA55_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA56_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA57_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA58_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA59_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA60_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA61_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA62_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA63_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA64_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA65_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA66_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA67_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA68_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA69_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA70_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA71_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA72_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA73_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA74_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA75_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA76_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA77_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA78_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA79_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA80_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA81_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA82_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA83_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA84_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA85_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA86_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA87_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA88_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA89_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA90_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA91_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA92_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA93_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA94_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA95_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA96_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA97_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA98_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA99_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA100_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA101_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA102_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA103_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA104_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA105_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA106_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA107_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA108_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA109_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA110_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA111_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA112_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA113_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA114_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA115_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA116_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA117_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA118_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA119_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA120_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA121_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA122_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA123_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA124_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA125_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA126_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDATA127_GlitchData : VitalGlitchDataType;
	variable  APUFCMLOADDVALID_GlitchData : VitalGlitchDataType;
	variable  APUFCMMSRFE0_GlitchData : VitalGlitchDataType;
	variable  APUFCMMSRFE1_GlitchData : VitalGlitchDataType;
	variable  APUFCMNEXTINSTRREADY_GlitchData : VitalGlitchDataType;
	variable  APUFCMOPERANDVALID_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA0_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA1_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA2_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA3_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA4_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA5_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA6_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA7_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA8_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA9_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA10_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA11_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA12_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA13_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA14_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA15_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA16_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA17_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA18_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA19_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA20_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA21_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA22_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA23_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA24_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA25_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA26_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA27_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA28_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA29_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA30_GlitchData : VitalGlitchDataType;
	variable  APUFCMRADATA31_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA0_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA1_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA2_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA3_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA4_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA5_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA6_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA7_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA8_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA9_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA10_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA11_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA12_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA13_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA14_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA15_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA16_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA17_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA18_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA19_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA20_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA21_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA22_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA23_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA24_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA25_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA26_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA27_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA28_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA29_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA30_GlitchData : VitalGlitchDataType;
	variable  APUFCMRBDATA31_GlitchData : VitalGlitchDataType;
	variable  APUFCMWRITEBACKOK_GlitchData : VitalGlitchDataType;
	variable  C440CPMCORESLEEPREQ_GlitchData : VitalGlitchDataType;
	variable  C440CPMDECIRPTREQ_GlitchData : VitalGlitchDataType;
	variable  C440CPMFITIRPTREQ_GlitchData : VitalGlitchDataType;
	variable  C440CPMMSRCE_GlitchData : VitalGlitchDataType;
	variable  C440CPMMSREE_GlitchData : VitalGlitchDataType;
	variable  C440CPMTIMERRESETREQ_GlitchData : VitalGlitchDataType;
	variable  C440CPMWDIRPTREQ_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL0_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL1_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL2_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL3_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL4_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL5_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL6_GlitchData : VitalGlitchDataType;
	variable  C440DBGSYSTEMCONTROL7_GlitchData : VitalGlitchDataType;
	variable  C440JTGTDO_GlitchData : VitalGlitchDataType;
	variable  C440JTGTDOEN_GlitchData : VitalGlitchDataType;
	variable  C440MACHINECHECK_GlitchData : VitalGlitchDataType;
	variable  C440RSTCHIPRESETREQ_GlitchData : VitalGlitchDataType;
	variable  C440RSTCORERESETREQ_GlitchData : VitalGlitchDataType;
	variable  C440RSTSYSTEMRESETREQ_GlitchData : VitalGlitchDataType;
	variable  C440TRCBRANCHSTATUS0_GlitchData : VitalGlitchDataType;
	variable  C440TRCBRANCHSTATUS1_GlitchData : VitalGlitchDataType;
	variable  C440TRCBRANCHSTATUS2_GlitchData : VitalGlitchDataType;
	variable  C440TRCCYCLE_GlitchData : VitalGlitchDataType;
	variable  C440TRCEXECUTIONSTATUS0_GlitchData : VitalGlitchDataType;
	variable  C440TRCEXECUTIONSTATUS1_GlitchData : VitalGlitchDataType;
	variable  C440TRCEXECUTIONSTATUS2_GlitchData : VitalGlitchDataType;
	variable  C440TRCEXECUTIONSTATUS3_GlitchData : VitalGlitchDataType;
	variable  C440TRCEXECUTIONSTATUS4_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRACESTATUS0_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRACESTATUS1_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRACESTATUS2_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRACESTATUS3_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRACESTATUS4_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRACESTATUS5_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRACESTATUS6_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTOUT_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE0_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE1_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE2_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE3_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE4_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE5_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE6_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE7_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE8_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE9_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE10_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE11_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE12_GlitchData : VitalGlitchDataType;
	variable  C440TRCTRIGGEREVENTTYPE13_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS0_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS1_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS2_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS3_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS4_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS5_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS6_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS7_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS8_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS9_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS10_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS11_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS12_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS13_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS14_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS15_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS16_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS17_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS18_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS19_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS20_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS21_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS22_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS23_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS24_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS25_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS26_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS27_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS28_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS29_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS30_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS31_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS32_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS33_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS34_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESS35_GlitchData : VitalGlitchDataType;
	variable  MIMCADDRESSVALID_GlitchData : VitalGlitchDataType;
	variable  MIMCBANKCONFLICT_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE0_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE1_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE2_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE3_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE4_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE5_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE6_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE7_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE8_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE9_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE10_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE11_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE12_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE13_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE14_GlitchData : VitalGlitchDataType;
	variable  MIMCBYTEENABLE15_GlitchData : VitalGlitchDataType;
	variable  MIMCREADNOTWRITE_GlitchData : VitalGlitchDataType;
	variable  MIMCROWCONFLICT_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA0_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA1_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA2_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA3_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA4_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA5_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA6_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA7_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA8_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA9_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA10_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA11_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA12_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA13_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA14_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA15_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA16_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA17_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA18_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA19_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA20_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA21_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA22_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA23_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA24_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA25_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA26_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA27_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA28_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA29_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA30_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA31_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA32_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA33_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA34_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA35_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA36_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA37_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA38_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA39_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA40_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA41_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA42_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA43_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA44_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA45_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA46_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA47_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA48_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA49_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA50_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA51_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA52_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA53_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA54_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA55_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA56_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA57_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA58_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA59_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA60_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA61_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA62_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA63_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA64_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA65_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA66_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA67_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA68_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA69_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA70_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA71_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA72_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA73_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA74_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA75_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA76_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA77_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA78_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA79_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA80_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA81_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA82_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA83_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA84_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA85_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA86_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA87_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA88_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA89_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA90_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA91_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA92_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA93_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA94_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA95_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA96_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA97_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA98_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA99_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA100_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA101_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA102_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA103_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA104_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA105_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA106_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA107_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA108_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA109_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA110_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA111_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA112_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA113_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA114_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA115_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA116_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA117_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA118_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA119_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA120_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA121_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA122_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA123_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA124_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA125_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA126_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATA127_GlitchData : VitalGlitchDataType;
	variable  MIMCWRITEDATAVALID_GlitchData : VitalGlitchDataType;
	variable  PPCCPMINTERCONNECTBUSY_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRACK_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRTIMEOUTWAIT_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN0_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN1_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN2_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN3_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN4_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN5_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN6_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN7_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN8_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN9_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN10_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN11_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN12_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN13_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN14_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN15_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN16_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN17_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN18_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN19_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN20_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN21_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN22_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN23_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN24_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN25_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN26_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN27_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN28_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN29_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN30_GlitchData : VitalGlitchDataType;
	variable  PPCDSDCRDBUSIN31_GlitchData : VitalGlitchDataType;
	variable  PPCEICINTERCONNECTIRQ_GlitchData : VitalGlitchDataType;
begin

     if (TimingChecksOn) then
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS0RNW_CPMPPCS0PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS0RNW_CPMPPCS0PLBCLK_posedge,
	TestSignal     => PLBPPCS0RNW,
	TestSignalName => "PLBPPCS0RNW",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName  => "CPMPPCS0PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS0RNW_CPMPPCS0PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS0RNW_CPMPPCS0PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS0RNW_CPMPPCS0PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS0RNW_CPMPPCS0PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS1RNW_CPMPPCS1PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS1RNW_CPMPPCS1PLBCLK_posedge,
	TestSignal     => PLBPPCS1RNW,
	TestSignalName => "PLBPPCS1RNW",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName  => "CPMPPCS1PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS1RNW_CPMPPCS1PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS1RNW_CPMPPCS1PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS1RNW_CPMPPCS1PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS1RNW_CPMPPCS1PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_CPMINTERCONNECTCLKNTO1_CPMINTERCONNECTCLK_posedge,
	TimingData     => Tmkr_CPMINTERCONNECTCLKNTO1_CPMINTERCONNECTCLK_posedge,
	TestSignal     => CPMINTERCONNECTCLKNTO1,
	TestSignalName => "CPMINTERCONNECTCLKNTO1",
	TestDelay      => 0 ps,
	RefSignal => CPMINTERCONNECTCLK_dly,
	RefSignalName  => "CPMINTERCONNECTCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_CPMINTERCONNECTCLKNTO1_CPMINTERCONNECTCLK_posedge_posedge,
	SetupLow       => tsetup_CPMINTERCONNECTCLKNTO1_CPMINTERCONNECTCLK_negedge_posedge,
	HoldLow        => thold_CPMINTERCONNECTCLKNTO1_CPMINTERCONNECTCLK_posedge_posedge,
	HoldHigh       => thold_CPMINTERCONNECTCLKNTO1_CPMINTERCONNECTCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_DCRPPCDMACK_CPMDCRCLK_posedge,
	TimingData     => Tmkr_DCRPPCDMACK_CPMDCRCLK_posedge,
	TestSignal     => DCRPPCDMACK,
	TestSignalName => "DCRPPCDMACK",
	TestDelay      => 0 ps,
	RefSignal => CPMDCRCLK_dly,
	RefSignalName  => "CPMDCRCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_DCRPPCDMACK_CPMDCRCLK_posedge_posedge,
	SetupLow       => tsetup_DCRPPCDMACK_CPMDCRCLK_negedge_posedge,
	HoldLow        => thold_DCRPPCDMACK_CPMDCRCLK_posedge_posedge,
	HoldHigh       => thold_DCRPPCDMACK_CPMDCRCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN0_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN0_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(0),
	TestSignalName => "DCRPPCDMDBUSIN(0)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(0),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(0),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(0),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(0),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN1_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN1_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(1),
	TestSignalName => "DCRPPCDMDBUSIN(1)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(1),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(1),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(1),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(1),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN2_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN2_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(2),
	TestSignalName => "DCRPPCDMDBUSIN(2)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(2),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(2),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(2),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(2),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN3_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN3_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(3),
	TestSignalName => "DCRPPCDMDBUSIN(3)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(3),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(3),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(3),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(3),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN4_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN4_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(4),
	TestSignalName => "DCRPPCDMDBUSIN(4)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(4),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(4),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(4),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(4),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN5_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN5_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(5),
	TestSignalName => "DCRPPCDMDBUSIN(5)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(5),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(5),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(5),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(5),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN6_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN6_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(6),
	TestSignalName => "DCRPPCDMDBUSIN(6)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(6),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(6),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(6),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(6),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN7_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN7_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(7),
	TestSignalName => "DCRPPCDMDBUSIN(7)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(7),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(7),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(7),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(7),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN8_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN8_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(8),
	TestSignalName => "DCRPPCDMDBUSIN(8)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(8),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(8),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(8),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(8),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN9_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN9_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(9),
	TestSignalName => "DCRPPCDMDBUSIN(9)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(9),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(9),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(9),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(9),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN10_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN10_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(10),
	TestSignalName => "DCRPPCDMDBUSIN(10)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(10),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(10),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(10),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(10),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN11_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN11_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(11),
	TestSignalName => "DCRPPCDMDBUSIN(11)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(11),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(11),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(11),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(11),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN12_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN12_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(12),
	TestSignalName => "DCRPPCDMDBUSIN(12)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(12),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(12),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(12),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(12),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN13_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN13_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(13),
	TestSignalName => "DCRPPCDMDBUSIN(13)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(13),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(13),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(13),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(13),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN14_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN14_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(14),
	TestSignalName => "DCRPPCDMDBUSIN(14)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(14),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(14),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(14),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(14),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN15_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN15_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(15),
	TestSignalName => "DCRPPCDMDBUSIN(15)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(15),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(15),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(15),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(15),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN16_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN16_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(16),
	TestSignalName => "DCRPPCDMDBUSIN(16)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(16),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(16),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(16),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(16),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(16),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN17_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN17_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(17),
	TestSignalName => "DCRPPCDMDBUSIN(17)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(17),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(17),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(17),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(17),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(17),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN18_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN18_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(18),
	TestSignalName => "DCRPPCDMDBUSIN(18)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(18),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(18),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(18),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(18),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(18),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN19_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN19_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(19),
	TestSignalName => "DCRPPCDMDBUSIN(19)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(19),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(19),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(19),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(19),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(19),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN20_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN20_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(20),
	TestSignalName => "DCRPPCDMDBUSIN(20)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(20),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(20),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(20),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(20),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(20),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN21_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN21_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(21),
	TestSignalName => "DCRPPCDMDBUSIN(21)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(21),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(21),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(21),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(21),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(21),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN22_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN22_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(22),
	TestSignalName => "DCRPPCDMDBUSIN(22)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(22),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(22),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(22),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(22),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(22),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN23_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN23_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(23),
	TestSignalName => "DCRPPCDMDBUSIN(23)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(23),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(23),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(23),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(23),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(23),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN24_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN24_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(24),
	TestSignalName => "DCRPPCDMDBUSIN(24)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(24),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(24),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(24),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(24),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(24),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN25_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN25_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(25),
	TestSignalName => "DCRPPCDMDBUSIN(25)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(25),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(25),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(25),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(25),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(25),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN26_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN26_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(26),
	TestSignalName => "DCRPPCDMDBUSIN(26)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(26),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(26),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(26),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(26),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(26),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN27_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN27_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(27),
	TestSignalName => "DCRPPCDMDBUSIN(27)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(27),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(27),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(27),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(27),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(27),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN28_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN28_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(28),
	TestSignalName => "DCRPPCDMDBUSIN(28)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(28),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(28),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(28),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(28),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN29_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN29_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(29),
	TestSignalName => "DCRPPCDMDBUSIN(29)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(29),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(29),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(29),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(29),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN30_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN30_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(30),
	TestSignalName => "DCRPPCDMDBUSIN(30)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(30),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(30),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(30),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(30),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDMDBUSIN31_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDMDBUSIN31_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDMDBUSIN_dly(31),
	TestSignalName => "DCRPPCDMDBUSIN(31)",
	TestDelay => tisd_DCRPPCDMDBUSIN_CPMDCRCLK(31),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(31),
	SetupLow => tsetup_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(31),
	HoldLow => thold_DCRPPCDMDBUSIN_CPMDCRCLK_posedge_posedge(31),
	HoldHigh => thold_DCRPPCDMDBUSIN_CPMDCRCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_DCRPPCDMTIMEOUTWAIT_CPMDCRCLK_posedge,
	TimingData     => Tmkr_DCRPPCDMTIMEOUTWAIT_CPMDCRCLK_posedge,
	TestSignal     => DCRPPCDMTIMEOUTWAIT,
	TestSignalName => "DCRPPCDMTIMEOUTWAIT",
	TestDelay      => 0 ps,
	RefSignal => CPMDCRCLK_dly,
	RefSignalName  => "CPMDCRCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_DCRPPCDMTIMEOUTWAIT_CPMDCRCLK_posedge_posedge,
	SetupLow       => tsetup_DCRPPCDMTIMEOUTWAIT_CPMDCRCLK_negedge_posedge,
	HoldLow        => thold_DCRPPCDMTIMEOUTWAIT_CPMDCRCLK_posedge_posedge,
	HoldHigh       => thold_DCRPPCDMTIMEOUTWAIT_CPMDCRCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA0RSTENGINEREQ_CPMDMA0LLCLK_posedge,
	TimingData     => Tmkr_LLDMA0RSTENGINEREQ_CPMDMA0LLCLK_posedge,
	TestSignal     => LLDMA0RSTENGINEREQ,
	TestSignalName => "LLDMA0RSTENGINEREQ",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName  => "CPMDMA0LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA0RSTENGINEREQ_CPMDMA0LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA0RSTENGINEREQ_CPMDMA0LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA0RSTENGINEREQ_CPMDMA0LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA0RSTENGINEREQ_CPMDMA0LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD0_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD0_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(0),
	TestSignalName => "LLDMA0RXD(0)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(0),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(0),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(0),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(0),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD1_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD1_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(1),
	TestSignalName => "LLDMA0RXD(1)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(1),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(1),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(1),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(1),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD2_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD2_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(2),
	TestSignalName => "LLDMA0RXD(2)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(2),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(2),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(2),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(2),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD3_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD3_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(3),
	TestSignalName => "LLDMA0RXD(3)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(3),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(3),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(3),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(3),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD4_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD4_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(4),
	TestSignalName => "LLDMA0RXD(4)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(4),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(4),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(4),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(4),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD5_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD5_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(5),
	TestSignalName => "LLDMA0RXD(5)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(5),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(5),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(5),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(5),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD6_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD6_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(6),
	TestSignalName => "LLDMA0RXD(6)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(6),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(6),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(6),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(6),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD7_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD7_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(7),
	TestSignalName => "LLDMA0RXD(7)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(7),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(7),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(7),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(7),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD8_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD8_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(8),
	TestSignalName => "LLDMA0RXD(8)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(8),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(8),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(8),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(8),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD9_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD9_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(9),
	TestSignalName => "LLDMA0RXD(9)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(9),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(9),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(9),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(9),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD10_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD10_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(10),
	TestSignalName => "LLDMA0RXD(10)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(10),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(10),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(10),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(10),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD11_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD11_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(11),
	TestSignalName => "LLDMA0RXD(11)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(11),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(11),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(11),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(11),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD12_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD12_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(12),
	TestSignalName => "LLDMA0RXD(12)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(12),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(12),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(12),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(12),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD13_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD13_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(13),
	TestSignalName => "LLDMA0RXD(13)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(13),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(13),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(13),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(13),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD14_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD14_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(14),
	TestSignalName => "LLDMA0RXD(14)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(14),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(14),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(14),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(14),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD15_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD15_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(15),
	TestSignalName => "LLDMA0RXD(15)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(15),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(15),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(15),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(15),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD16_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD16_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(16),
	TestSignalName => "LLDMA0RXD(16)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(16),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(16),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(16),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(16),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(16),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD17_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD17_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(17),
	TestSignalName => "LLDMA0RXD(17)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(17),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(17),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(17),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(17),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(17),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD18_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD18_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(18),
	TestSignalName => "LLDMA0RXD(18)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(18),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(18),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(18),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(18),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(18),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD19_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD19_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(19),
	TestSignalName => "LLDMA0RXD(19)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(19),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(19),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(19),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(19),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(19),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD20_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD20_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(20),
	TestSignalName => "LLDMA0RXD(20)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(20),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(20),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(20),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(20),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(20),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD21_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD21_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(21),
	TestSignalName => "LLDMA0RXD(21)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(21),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(21),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(21),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(21),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(21),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD22_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD22_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(22),
	TestSignalName => "LLDMA0RXD(22)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(22),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(22),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(22),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(22),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(22),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD23_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD23_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(23),
	TestSignalName => "LLDMA0RXD(23)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(23),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(23),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(23),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(23),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(23),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD24_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD24_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(24),
	TestSignalName => "LLDMA0RXD(24)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(24),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(24),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(24),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(24),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(24),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD25_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD25_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(25),
	TestSignalName => "LLDMA0RXD(25)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(25),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(25),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(25),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(25),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(25),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD26_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD26_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(26),
	TestSignalName => "LLDMA0RXD(26)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(26),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(26),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(26),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(26),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(26),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD27_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD27_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(27),
	TestSignalName => "LLDMA0RXD(27)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(27),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(27),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(27),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(27),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(27),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD28_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD28_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(28),
	TestSignalName => "LLDMA0RXD(28)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(28),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(28),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(28),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(28),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD29_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD29_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(29),
	TestSignalName => "LLDMA0RXD(29)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(29),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(29),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(29),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(29),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD30_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD30_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(30),
	TestSignalName => "LLDMA0RXD(30)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(30),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(30),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(30),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(30),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXD31_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXD31_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXD_dly(31),
	TestSignalName => "LLDMA0RXD(31)",
	TestDelay => tisd_LLDMA0RXD_CPMDMA0LLCLK(31),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(31),
	SetupLow => tsetup_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(31),
	HoldLow => thold_LLDMA0RXD_CPMDMA0LLCLK_posedge_posedge(31),
	HoldHigh => thold_LLDMA0RXD_CPMDMA0LLCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA0RXEOFN_CPMDMA0LLCLK_posedge,
	TimingData     => Tmkr_LLDMA0RXEOFN_CPMDMA0LLCLK_posedge,
	TestSignal     => LLDMA0RXEOFN,
	TestSignalName => "LLDMA0RXEOFN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName  => "CPMDMA0LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA0RXEOFN_CPMDMA0LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA0RXEOFN_CPMDMA0LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA0RXEOFN_CPMDMA0LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA0RXEOFN_CPMDMA0LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA0RXEOPN_CPMDMA0LLCLK_posedge,
	TimingData     => Tmkr_LLDMA0RXEOPN_CPMDMA0LLCLK_posedge,
	TestSignal     => LLDMA0RXEOPN,
	TestSignalName => "LLDMA0RXEOPN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName  => "CPMDMA0LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA0RXEOPN_CPMDMA0LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA0RXEOPN_CPMDMA0LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA0RXEOPN_CPMDMA0LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA0RXEOPN_CPMDMA0LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXREM0_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXREM0_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXREM_dly(0),
	TestSignalName => "LLDMA0RXREM(0)",
	TestDelay => tisd_LLDMA0RXREM_CPMDMA0LLCLK(0),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXREM_CPMDMA0LLCLK_posedge_posedge(0),
	SetupLow => tsetup_LLDMA0RXREM_CPMDMA0LLCLK_negedge_posedge(0),
	HoldLow => thold_LLDMA0RXREM_CPMDMA0LLCLK_posedge_posedge(0),
	HoldHigh => thold_LLDMA0RXREM_CPMDMA0LLCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXREM1_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXREM1_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXREM_dly(1),
	TestSignalName => "LLDMA0RXREM(1)",
	TestDelay => tisd_LLDMA0RXREM_CPMDMA0LLCLK(1),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXREM_CPMDMA0LLCLK_posedge_posedge(1),
	SetupLow => tsetup_LLDMA0RXREM_CPMDMA0LLCLK_negedge_posedge(1),
	HoldLow => thold_LLDMA0RXREM_CPMDMA0LLCLK_posedge_posedge(1),
	HoldHigh => thold_LLDMA0RXREM_CPMDMA0LLCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXREM2_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXREM2_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXREM_dly(2),
	TestSignalName => "LLDMA0RXREM(2)",
	TestDelay => tisd_LLDMA0RXREM_CPMDMA0LLCLK(2),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXREM_CPMDMA0LLCLK_posedge_posedge(2),
	SetupLow => tsetup_LLDMA0RXREM_CPMDMA0LLCLK_negedge_posedge(2),
	HoldLow => thold_LLDMA0RXREM_CPMDMA0LLCLK_posedge_posedge(2),
	HoldHigh => thold_LLDMA0RXREM_CPMDMA0LLCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA0RXREM3_CPMDMA0LLCLK_posedge,
	TimingData => Tmkr_LLDMA0RXREM3_CPMDMA0LLCLK_posedge,
	TestSignal => LLDMA0RXREM_dly(3),
	TestSignalName => "LLDMA0RXREM(3)",
	TestDelay => tisd_LLDMA0RXREM_CPMDMA0LLCLK(3),
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName => "CPMDMA0LLCLK",
	RefDelay => ticd_CPMDMA0LLCLK,
	SetupHigh => tsetup_LLDMA0RXREM_CPMDMA0LLCLK_posedge_posedge(3),
	SetupLow => tsetup_LLDMA0RXREM_CPMDMA0LLCLK_negedge_posedge(3),
	HoldLow => thold_LLDMA0RXREM_CPMDMA0LLCLK_posedge_posedge(3),
	HoldHigh => thold_LLDMA0RXREM_CPMDMA0LLCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA0RXSOFN_CPMDMA0LLCLK_posedge,
	TimingData     => Tmkr_LLDMA0RXSOFN_CPMDMA0LLCLK_posedge,
	TestSignal     => LLDMA0RXSOFN,
	TestSignalName => "LLDMA0RXSOFN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName  => "CPMDMA0LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA0RXSOFN_CPMDMA0LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA0RXSOFN_CPMDMA0LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA0RXSOFN_CPMDMA0LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA0RXSOFN_CPMDMA0LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA0RXSOPN_CPMDMA0LLCLK_posedge,
	TimingData     => Tmkr_LLDMA0RXSOPN_CPMDMA0LLCLK_posedge,
	TestSignal     => LLDMA0RXSOPN,
	TestSignalName => "LLDMA0RXSOPN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName  => "CPMDMA0LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA0RXSOPN_CPMDMA0LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA0RXSOPN_CPMDMA0LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA0RXSOPN_CPMDMA0LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA0RXSOPN_CPMDMA0LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA0RXSRCRDYN_CPMDMA0LLCLK_posedge,
	TimingData     => Tmkr_LLDMA0RXSRCRDYN_CPMDMA0LLCLK_posedge,
	TestSignal     => LLDMA0RXSRCRDYN,
	TestSignalName => "LLDMA0RXSRCRDYN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName  => "CPMDMA0LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA0RXSRCRDYN_CPMDMA0LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA0RXSRCRDYN_CPMDMA0LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA0RXSRCRDYN_CPMDMA0LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA0RXSRCRDYN_CPMDMA0LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA0TXDSTRDYN_CPMDMA0LLCLK_posedge,
	TimingData     => Tmkr_LLDMA0TXDSTRDYN_CPMDMA0LLCLK_posedge,
	TestSignal     => LLDMA0TXDSTRDYN,
	TestSignalName => "LLDMA0TXDSTRDYN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA0LLCLK_dly,
	RefSignalName  => "CPMDMA0LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA0TXDSTRDYN_CPMDMA0LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA0TXDSTRDYN_CPMDMA0LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA0TXDSTRDYN_CPMDMA0LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA0TXDSTRDYN_CPMDMA0LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA1RSTENGINEREQ_CPMDMA1LLCLK_posedge,
	TimingData     => Tmkr_LLDMA1RSTENGINEREQ_CPMDMA1LLCLK_posedge,
	TestSignal     => LLDMA1RSTENGINEREQ,
	TestSignalName => "LLDMA1RSTENGINEREQ",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName  => "CPMDMA1LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA1RSTENGINEREQ_CPMDMA1LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA1RSTENGINEREQ_CPMDMA1LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA1RSTENGINEREQ_CPMDMA1LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA1RSTENGINEREQ_CPMDMA1LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD0_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD0_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(0),
	TestSignalName => "LLDMA1RXD(0)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(0),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(0),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(0),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(0),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD1_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD1_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(1),
	TestSignalName => "LLDMA1RXD(1)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(1),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(1),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(1),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(1),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD2_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD2_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(2),
	TestSignalName => "LLDMA1RXD(2)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(2),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(2),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(2),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(2),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD3_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD3_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(3),
	TestSignalName => "LLDMA1RXD(3)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(3),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(3),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(3),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(3),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD4_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD4_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(4),
	TestSignalName => "LLDMA1RXD(4)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(4),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(4),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(4),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(4),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD5_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD5_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(5),
	TestSignalName => "LLDMA1RXD(5)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(5),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(5),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(5),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(5),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD6_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD6_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(6),
	TestSignalName => "LLDMA1RXD(6)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(6),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(6),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(6),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(6),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD7_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD7_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(7),
	TestSignalName => "LLDMA1RXD(7)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(7),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(7),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(7),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(7),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD8_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD8_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(8),
	TestSignalName => "LLDMA1RXD(8)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(8),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(8),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(8),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(8),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD9_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD9_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(9),
	TestSignalName => "LLDMA1RXD(9)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(9),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(9),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(9),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(9),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD10_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD10_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(10),
	TestSignalName => "LLDMA1RXD(10)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(10),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(10),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(10),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(10),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD11_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD11_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(11),
	TestSignalName => "LLDMA1RXD(11)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(11),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(11),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(11),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(11),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD12_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD12_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(12),
	TestSignalName => "LLDMA1RXD(12)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(12),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(12),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(12),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(12),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD13_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD13_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(13),
	TestSignalName => "LLDMA1RXD(13)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(13),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(13),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(13),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(13),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD14_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD14_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(14),
	TestSignalName => "LLDMA1RXD(14)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(14),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(14),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(14),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(14),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD15_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD15_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(15),
	TestSignalName => "LLDMA1RXD(15)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(15),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(15),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(15),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(15),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD16_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD16_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(16),
	TestSignalName => "LLDMA1RXD(16)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(16),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(16),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(16),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(16),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(16),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD17_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD17_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(17),
	TestSignalName => "LLDMA1RXD(17)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(17),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(17),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(17),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(17),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(17),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD18_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD18_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(18),
	TestSignalName => "LLDMA1RXD(18)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(18),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(18),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(18),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(18),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(18),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD19_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD19_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(19),
	TestSignalName => "LLDMA1RXD(19)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(19),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(19),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(19),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(19),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(19),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD20_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD20_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(20),
	TestSignalName => "LLDMA1RXD(20)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(20),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(20),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(20),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(20),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(20),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD21_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD21_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(21),
	TestSignalName => "LLDMA1RXD(21)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(21),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(21),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(21),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(21),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(21),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD22_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD22_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(22),
	TestSignalName => "LLDMA1RXD(22)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(22),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(22),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(22),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(22),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(22),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD23_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD23_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(23),
	TestSignalName => "LLDMA1RXD(23)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(23),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(23),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(23),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(23),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(23),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD24_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD24_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(24),
	TestSignalName => "LLDMA1RXD(24)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(24),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(24),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(24),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(24),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(24),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD25_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD25_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(25),
	TestSignalName => "LLDMA1RXD(25)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(25),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(25),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(25),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(25),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(25),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD26_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD26_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(26),
	TestSignalName => "LLDMA1RXD(26)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(26),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(26),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(26),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(26),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(26),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD27_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD27_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(27),
	TestSignalName => "LLDMA1RXD(27)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(27),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(27),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(27),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(27),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(27),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD28_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD28_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(28),
	TestSignalName => "LLDMA1RXD(28)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(28),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(28),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(28),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(28),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD29_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD29_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(29),
	TestSignalName => "LLDMA1RXD(29)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(29),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(29),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(29),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(29),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD30_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD30_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(30),
	TestSignalName => "LLDMA1RXD(30)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(30),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(30),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(30),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(30),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXD31_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXD31_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXD_dly(31),
	TestSignalName => "LLDMA1RXD(31)",
	TestDelay => tisd_LLDMA1RXD_CPMDMA1LLCLK(31),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(31),
	SetupLow => tsetup_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(31),
	HoldLow => thold_LLDMA1RXD_CPMDMA1LLCLK_posedge_posedge(31),
	HoldHigh => thold_LLDMA1RXD_CPMDMA1LLCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA1RXEOFN_CPMDMA1LLCLK_posedge,
	TimingData     => Tmkr_LLDMA1RXEOFN_CPMDMA1LLCLK_posedge,
	TestSignal     => LLDMA1RXEOFN,
	TestSignalName => "LLDMA1RXEOFN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName  => "CPMDMA1LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA1RXEOFN_CPMDMA1LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA1RXEOFN_CPMDMA1LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA1RXEOFN_CPMDMA1LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA1RXEOFN_CPMDMA1LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA1RXEOPN_CPMDMA1LLCLK_posedge,
	TimingData     => Tmkr_LLDMA1RXEOPN_CPMDMA1LLCLK_posedge,
	TestSignal     => LLDMA1RXEOPN,
	TestSignalName => "LLDMA1RXEOPN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName  => "CPMDMA1LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA1RXEOPN_CPMDMA1LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA1RXEOPN_CPMDMA1LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA1RXEOPN_CPMDMA1LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA1RXEOPN_CPMDMA1LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXREM0_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXREM0_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXREM_dly(0),
	TestSignalName => "LLDMA1RXREM(0)",
	TestDelay => tisd_LLDMA1RXREM_CPMDMA1LLCLK(0),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXREM_CPMDMA1LLCLK_posedge_posedge(0),
	SetupLow => tsetup_LLDMA1RXREM_CPMDMA1LLCLK_negedge_posedge(0),
	HoldLow => thold_LLDMA1RXREM_CPMDMA1LLCLK_posedge_posedge(0),
	HoldHigh => thold_LLDMA1RXREM_CPMDMA1LLCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXREM1_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXREM1_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXREM_dly(1),
	TestSignalName => "LLDMA1RXREM(1)",
	TestDelay => tisd_LLDMA1RXREM_CPMDMA1LLCLK(1),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXREM_CPMDMA1LLCLK_posedge_posedge(1),
	SetupLow => tsetup_LLDMA1RXREM_CPMDMA1LLCLK_negedge_posedge(1),
	HoldLow => thold_LLDMA1RXREM_CPMDMA1LLCLK_posedge_posedge(1),
	HoldHigh => thold_LLDMA1RXREM_CPMDMA1LLCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXREM2_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXREM2_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXREM_dly(2),
	TestSignalName => "LLDMA1RXREM(2)",
	TestDelay => tisd_LLDMA1RXREM_CPMDMA1LLCLK(2),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXREM_CPMDMA1LLCLK_posedge_posedge(2),
	SetupLow => tsetup_LLDMA1RXREM_CPMDMA1LLCLK_negedge_posedge(2),
	HoldLow => thold_LLDMA1RXREM_CPMDMA1LLCLK_posedge_posedge(2),
	HoldHigh => thold_LLDMA1RXREM_CPMDMA1LLCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA1RXREM3_CPMDMA1LLCLK_posedge,
	TimingData => Tmkr_LLDMA1RXREM3_CPMDMA1LLCLK_posedge,
	TestSignal => LLDMA1RXREM_dly(3),
	TestSignalName => "LLDMA1RXREM(3)",
	TestDelay => tisd_LLDMA1RXREM_CPMDMA1LLCLK(3),
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName => "CPMDMA1LLCLK",
	RefDelay => ticd_CPMDMA1LLCLK,
	SetupHigh => tsetup_LLDMA1RXREM_CPMDMA1LLCLK_posedge_posedge(3),
	SetupLow => tsetup_LLDMA1RXREM_CPMDMA1LLCLK_negedge_posedge(3),
	HoldLow => thold_LLDMA1RXREM_CPMDMA1LLCLK_posedge_posedge(3),
	HoldHigh => thold_LLDMA1RXREM_CPMDMA1LLCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA1RXSOFN_CPMDMA1LLCLK_posedge,
	TimingData     => Tmkr_LLDMA1RXSOFN_CPMDMA1LLCLK_posedge,
	TestSignal     => LLDMA1RXSOFN,
	TestSignalName => "LLDMA1RXSOFN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName  => "CPMDMA1LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA1RXSOFN_CPMDMA1LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA1RXSOFN_CPMDMA1LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA1RXSOFN_CPMDMA1LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA1RXSOFN_CPMDMA1LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA1RXSOPN_CPMDMA1LLCLK_posedge,
	TimingData     => Tmkr_LLDMA1RXSOPN_CPMDMA1LLCLK_posedge,
	TestSignal     => LLDMA1RXSOPN,
	TestSignalName => "LLDMA1RXSOPN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName  => "CPMDMA1LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA1RXSOPN_CPMDMA1LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA1RXSOPN_CPMDMA1LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA1RXSOPN_CPMDMA1LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA1RXSOPN_CPMDMA1LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA1RXSRCRDYN_CPMDMA1LLCLK_posedge,
	TimingData     => Tmkr_LLDMA1RXSRCRDYN_CPMDMA1LLCLK_posedge,
	TestSignal     => LLDMA1RXSRCRDYN,
	TestSignalName => "LLDMA1RXSRCRDYN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName  => "CPMDMA1LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA1RXSRCRDYN_CPMDMA1LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA1RXSRCRDYN_CPMDMA1LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA1RXSRCRDYN_CPMDMA1LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA1RXSRCRDYN_CPMDMA1LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA1TXDSTRDYN_CPMDMA1LLCLK_posedge,
	TimingData     => Tmkr_LLDMA1TXDSTRDYN_CPMDMA1LLCLK_posedge,
	TestSignal     => LLDMA1TXDSTRDYN,
	TestSignalName => "LLDMA1TXDSTRDYN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA1LLCLK_dly,
	RefSignalName  => "CPMDMA1LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA1TXDSTRDYN_CPMDMA1LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA1TXDSTRDYN_CPMDMA1LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA1TXDSTRDYN_CPMDMA1LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA1TXDSTRDYN_CPMDMA1LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA2RSTENGINEREQ_CPMDMA2LLCLK_posedge,
	TimingData     => Tmkr_LLDMA2RSTENGINEREQ_CPMDMA2LLCLK_posedge,
	TestSignal     => LLDMA2RSTENGINEREQ,
	TestSignalName => "LLDMA2RSTENGINEREQ",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName  => "CPMDMA2LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA2RSTENGINEREQ_CPMDMA2LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA2RSTENGINEREQ_CPMDMA2LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA2RSTENGINEREQ_CPMDMA2LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA2RSTENGINEREQ_CPMDMA2LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD0_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD0_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(0),
	TestSignalName => "LLDMA2RXD(0)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(0),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(0),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(0),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(0),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD1_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD1_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(1),
	TestSignalName => "LLDMA2RXD(1)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(1),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(1),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(1),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(1),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD2_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD2_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(2),
	TestSignalName => "LLDMA2RXD(2)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(2),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(2),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(2),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(2),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD3_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD3_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(3),
	TestSignalName => "LLDMA2RXD(3)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(3),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(3),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(3),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(3),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD4_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD4_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(4),
	TestSignalName => "LLDMA2RXD(4)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(4),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(4),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(4),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(4),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD5_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD5_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(5),
	TestSignalName => "LLDMA2RXD(5)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(5),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(5),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(5),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(5),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD6_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD6_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(6),
	TestSignalName => "LLDMA2RXD(6)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(6),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(6),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(6),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(6),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD7_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD7_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(7),
	TestSignalName => "LLDMA2RXD(7)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(7),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(7),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(7),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(7),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD8_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD8_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(8),
	TestSignalName => "LLDMA2RXD(8)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(8),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(8),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(8),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(8),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD9_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD9_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(9),
	TestSignalName => "LLDMA2RXD(9)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(9),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(9),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(9),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(9),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD10_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD10_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(10),
	TestSignalName => "LLDMA2RXD(10)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(10),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(10),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(10),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(10),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD11_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD11_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(11),
	TestSignalName => "LLDMA2RXD(11)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(11),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(11),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(11),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(11),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD12_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD12_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(12),
	TestSignalName => "LLDMA2RXD(12)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(12),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(12),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(12),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(12),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD13_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD13_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(13),
	TestSignalName => "LLDMA2RXD(13)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(13),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(13),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(13),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(13),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD14_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD14_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(14),
	TestSignalName => "LLDMA2RXD(14)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(14),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(14),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(14),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(14),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD15_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD15_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(15),
	TestSignalName => "LLDMA2RXD(15)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(15),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(15),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(15),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(15),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD16_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD16_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(16),
	TestSignalName => "LLDMA2RXD(16)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(16),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(16),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(16),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(16),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(16),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD17_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD17_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(17),
	TestSignalName => "LLDMA2RXD(17)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(17),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(17),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(17),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(17),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(17),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD18_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD18_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(18),
	TestSignalName => "LLDMA2RXD(18)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(18),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(18),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(18),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(18),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(18),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD19_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD19_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(19),
	TestSignalName => "LLDMA2RXD(19)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(19),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(19),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(19),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(19),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(19),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD20_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD20_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(20),
	TestSignalName => "LLDMA2RXD(20)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(20),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(20),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(20),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(20),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(20),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD21_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD21_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(21),
	TestSignalName => "LLDMA2RXD(21)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(21),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(21),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(21),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(21),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(21),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD22_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD22_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(22),
	TestSignalName => "LLDMA2RXD(22)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(22),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(22),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(22),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(22),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(22),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD23_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD23_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(23),
	TestSignalName => "LLDMA2RXD(23)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(23),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(23),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(23),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(23),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(23),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD24_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD24_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(24),
	TestSignalName => "LLDMA2RXD(24)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(24),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(24),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(24),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(24),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(24),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD25_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD25_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(25),
	TestSignalName => "LLDMA2RXD(25)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(25),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(25),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(25),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(25),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(25),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD26_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD26_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(26),
	TestSignalName => "LLDMA2RXD(26)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(26),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(26),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(26),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(26),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(26),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD27_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD27_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(27),
	TestSignalName => "LLDMA2RXD(27)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(27),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(27),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(27),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(27),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(27),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD28_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD28_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(28),
	TestSignalName => "LLDMA2RXD(28)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(28),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(28),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(28),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(28),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD29_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD29_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(29),
	TestSignalName => "LLDMA2RXD(29)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(29),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(29),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(29),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(29),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD30_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD30_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(30),
	TestSignalName => "LLDMA2RXD(30)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(30),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(30),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(30),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(30),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXD31_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXD31_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXD_dly(31),
	TestSignalName => "LLDMA2RXD(31)",
	TestDelay => tisd_LLDMA2RXD_CPMDMA2LLCLK(31),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(31),
	SetupLow => tsetup_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(31),
	HoldLow => thold_LLDMA2RXD_CPMDMA2LLCLK_posedge_posedge(31),
	HoldHigh => thold_LLDMA2RXD_CPMDMA2LLCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA2RXEOFN_CPMDMA2LLCLK_posedge,
	TimingData     => Tmkr_LLDMA2RXEOFN_CPMDMA2LLCLK_posedge,
	TestSignal     => LLDMA2RXEOFN,
	TestSignalName => "LLDMA2RXEOFN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName  => "CPMDMA2LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA2RXEOFN_CPMDMA2LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA2RXEOFN_CPMDMA2LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA2RXEOFN_CPMDMA2LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA2RXEOFN_CPMDMA2LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA2RXEOPN_CPMDMA2LLCLK_posedge,
	TimingData     => Tmkr_LLDMA2RXEOPN_CPMDMA2LLCLK_posedge,
	TestSignal     => LLDMA2RXEOPN,
	TestSignalName => "LLDMA2RXEOPN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName  => "CPMDMA2LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA2RXEOPN_CPMDMA2LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA2RXEOPN_CPMDMA2LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA2RXEOPN_CPMDMA2LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA2RXEOPN_CPMDMA2LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXREM0_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXREM0_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXREM_dly(0),
	TestSignalName => "LLDMA2RXREM(0)",
	TestDelay => tisd_LLDMA2RXREM_CPMDMA2LLCLK(0),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXREM_CPMDMA2LLCLK_posedge_posedge(0),
	SetupLow => tsetup_LLDMA2RXREM_CPMDMA2LLCLK_negedge_posedge(0),
	HoldLow => thold_LLDMA2RXREM_CPMDMA2LLCLK_posedge_posedge(0),
	HoldHigh => thold_LLDMA2RXREM_CPMDMA2LLCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXREM1_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXREM1_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXREM_dly(1),
	TestSignalName => "LLDMA2RXREM(1)",
	TestDelay => tisd_LLDMA2RXREM_CPMDMA2LLCLK(1),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXREM_CPMDMA2LLCLK_posedge_posedge(1),
	SetupLow => tsetup_LLDMA2RXREM_CPMDMA2LLCLK_negedge_posedge(1),
	HoldLow => thold_LLDMA2RXREM_CPMDMA2LLCLK_posedge_posedge(1),
	HoldHigh => thold_LLDMA2RXREM_CPMDMA2LLCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXREM2_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXREM2_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXREM_dly(2),
	TestSignalName => "LLDMA2RXREM(2)",
	TestDelay => tisd_LLDMA2RXREM_CPMDMA2LLCLK(2),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXREM_CPMDMA2LLCLK_posedge_posedge(2),
	SetupLow => tsetup_LLDMA2RXREM_CPMDMA2LLCLK_negedge_posedge(2),
	HoldLow => thold_LLDMA2RXREM_CPMDMA2LLCLK_posedge_posedge(2),
	HoldHigh => thold_LLDMA2RXREM_CPMDMA2LLCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA2RXREM3_CPMDMA2LLCLK_posedge,
	TimingData => Tmkr_LLDMA2RXREM3_CPMDMA2LLCLK_posedge,
	TestSignal => LLDMA2RXREM_dly(3),
	TestSignalName => "LLDMA2RXREM(3)",
	TestDelay => tisd_LLDMA2RXREM_CPMDMA2LLCLK(3),
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName => "CPMDMA2LLCLK",
	RefDelay => ticd_CPMDMA2LLCLK,
	SetupHigh => tsetup_LLDMA2RXREM_CPMDMA2LLCLK_posedge_posedge(3),
	SetupLow => tsetup_LLDMA2RXREM_CPMDMA2LLCLK_negedge_posedge(3),
	HoldLow => thold_LLDMA2RXREM_CPMDMA2LLCLK_posedge_posedge(3),
	HoldHigh => thold_LLDMA2RXREM_CPMDMA2LLCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA2RXSOFN_CPMDMA2LLCLK_posedge,
	TimingData     => Tmkr_LLDMA2RXSOFN_CPMDMA2LLCLK_posedge,
	TestSignal     => LLDMA2RXSOFN,
	TestSignalName => "LLDMA2RXSOFN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName  => "CPMDMA2LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA2RXSOFN_CPMDMA2LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA2RXSOFN_CPMDMA2LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA2RXSOFN_CPMDMA2LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA2RXSOFN_CPMDMA2LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA2RXSOPN_CPMDMA2LLCLK_posedge,
	TimingData     => Tmkr_LLDMA2RXSOPN_CPMDMA2LLCLK_posedge,
	TestSignal     => LLDMA2RXSOPN,
	TestSignalName => "LLDMA2RXSOPN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName  => "CPMDMA2LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA2RXSOPN_CPMDMA2LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA2RXSOPN_CPMDMA2LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA2RXSOPN_CPMDMA2LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA2RXSOPN_CPMDMA2LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA2RXSRCRDYN_CPMDMA2LLCLK_posedge,
	TimingData     => Tmkr_LLDMA2RXSRCRDYN_CPMDMA2LLCLK_posedge,
	TestSignal     => LLDMA2RXSRCRDYN,
	TestSignalName => "LLDMA2RXSRCRDYN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName  => "CPMDMA2LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA2RXSRCRDYN_CPMDMA2LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA2RXSRCRDYN_CPMDMA2LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA2RXSRCRDYN_CPMDMA2LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA2RXSRCRDYN_CPMDMA2LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA2TXDSTRDYN_CPMDMA2LLCLK_posedge,
	TimingData     => Tmkr_LLDMA2TXDSTRDYN_CPMDMA2LLCLK_posedge,
	TestSignal     => LLDMA2TXDSTRDYN,
	TestSignalName => "LLDMA2TXDSTRDYN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA2LLCLK_dly,
	RefSignalName  => "CPMDMA2LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA2TXDSTRDYN_CPMDMA2LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA2TXDSTRDYN_CPMDMA2LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA2TXDSTRDYN_CPMDMA2LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA2TXDSTRDYN_CPMDMA2LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA3RSTENGINEREQ_CPMDMA3LLCLK_posedge,
	TimingData     => Tmkr_LLDMA3RSTENGINEREQ_CPMDMA3LLCLK_posedge,
	TestSignal     => LLDMA3RSTENGINEREQ,
	TestSignalName => "LLDMA3RSTENGINEREQ",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName  => "CPMDMA3LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA3RSTENGINEREQ_CPMDMA3LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA3RSTENGINEREQ_CPMDMA3LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA3RSTENGINEREQ_CPMDMA3LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA3RSTENGINEREQ_CPMDMA3LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD0_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD0_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(0),
	TestSignalName => "LLDMA3RXD(0)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(0),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(0),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(0),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(0),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD1_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD1_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(1),
	TestSignalName => "LLDMA3RXD(1)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(1),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(1),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(1),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(1),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD2_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD2_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(2),
	TestSignalName => "LLDMA3RXD(2)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(2),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(2),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(2),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(2),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD3_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD3_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(3),
	TestSignalName => "LLDMA3RXD(3)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(3),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(3),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(3),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(3),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD4_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD4_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(4),
	TestSignalName => "LLDMA3RXD(4)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(4),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(4),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(4),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(4),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD5_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD5_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(5),
	TestSignalName => "LLDMA3RXD(5)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(5),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(5),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(5),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(5),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD6_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD6_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(6),
	TestSignalName => "LLDMA3RXD(6)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(6),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(6),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(6),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(6),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD7_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD7_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(7),
	TestSignalName => "LLDMA3RXD(7)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(7),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(7),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(7),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(7),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD8_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD8_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(8),
	TestSignalName => "LLDMA3RXD(8)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(8),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(8),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(8),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(8),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD9_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD9_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(9),
	TestSignalName => "LLDMA3RXD(9)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(9),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(9),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(9),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(9),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD10_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD10_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(10),
	TestSignalName => "LLDMA3RXD(10)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(10),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(10),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(10),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(10),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD11_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD11_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(11),
	TestSignalName => "LLDMA3RXD(11)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(11),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(11),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(11),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(11),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD12_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD12_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(12),
	TestSignalName => "LLDMA3RXD(12)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(12),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(12),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(12),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(12),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD13_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD13_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(13),
	TestSignalName => "LLDMA3RXD(13)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(13),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(13),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(13),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(13),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD14_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD14_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(14),
	TestSignalName => "LLDMA3RXD(14)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(14),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(14),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(14),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(14),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD15_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD15_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(15),
	TestSignalName => "LLDMA3RXD(15)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(15),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(15),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(15),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(15),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD16_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD16_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(16),
	TestSignalName => "LLDMA3RXD(16)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(16),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(16),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(16),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(16),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(16),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD17_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD17_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(17),
	TestSignalName => "LLDMA3RXD(17)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(17),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(17),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(17),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(17),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(17),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD18_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD18_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(18),
	TestSignalName => "LLDMA3RXD(18)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(18),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(18),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(18),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(18),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(18),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD19_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD19_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(19),
	TestSignalName => "LLDMA3RXD(19)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(19),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(19),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(19),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(19),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(19),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD20_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD20_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(20),
	TestSignalName => "LLDMA3RXD(20)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(20),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(20),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(20),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(20),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(20),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD21_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD21_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(21),
	TestSignalName => "LLDMA3RXD(21)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(21),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(21),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(21),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(21),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(21),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD22_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD22_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(22),
	TestSignalName => "LLDMA3RXD(22)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(22),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(22),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(22),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(22),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(22),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD23_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD23_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(23),
	TestSignalName => "LLDMA3RXD(23)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(23),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(23),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(23),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(23),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(23),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD24_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD24_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(24),
	TestSignalName => "LLDMA3RXD(24)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(24),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(24),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(24),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(24),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(24),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD25_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD25_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(25),
	TestSignalName => "LLDMA3RXD(25)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(25),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(25),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(25),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(25),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(25),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD26_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD26_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(26),
	TestSignalName => "LLDMA3RXD(26)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(26),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(26),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(26),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(26),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(26),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD27_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD27_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(27),
	TestSignalName => "LLDMA3RXD(27)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(27),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(27),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(27),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(27),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(27),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD28_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD28_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(28),
	TestSignalName => "LLDMA3RXD(28)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(28),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(28),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(28),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(28),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD29_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD29_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(29),
	TestSignalName => "LLDMA3RXD(29)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(29),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(29),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(29),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(29),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD30_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD30_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(30),
	TestSignalName => "LLDMA3RXD(30)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(30),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(30),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(30),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(30),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXD31_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXD31_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXD_dly(31),
	TestSignalName => "LLDMA3RXD(31)",
	TestDelay => tisd_LLDMA3RXD_CPMDMA3LLCLK(31),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(31),
	SetupLow => tsetup_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(31),
	HoldLow => thold_LLDMA3RXD_CPMDMA3LLCLK_posedge_posedge(31),
	HoldHigh => thold_LLDMA3RXD_CPMDMA3LLCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA3RXEOFN_CPMDMA3LLCLK_posedge,
	TimingData     => Tmkr_LLDMA3RXEOFN_CPMDMA3LLCLK_posedge,
	TestSignal     => LLDMA3RXEOFN,
	TestSignalName => "LLDMA3RXEOFN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName  => "CPMDMA3LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA3RXEOFN_CPMDMA3LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA3RXEOFN_CPMDMA3LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA3RXEOFN_CPMDMA3LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA3RXEOFN_CPMDMA3LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA3RXEOPN_CPMDMA3LLCLK_posedge,
	TimingData     => Tmkr_LLDMA3RXEOPN_CPMDMA3LLCLK_posedge,
	TestSignal     => LLDMA3RXEOPN,
	TestSignalName => "LLDMA3RXEOPN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName  => "CPMDMA3LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA3RXEOPN_CPMDMA3LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA3RXEOPN_CPMDMA3LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA3RXEOPN_CPMDMA3LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA3RXEOPN_CPMDMA3LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXREM0_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXREM0_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXREM_dly(0),
	TestSignalName => "LLDMA3RXREM(0)",
	TestDelay => tisd_LLDMA3RXREM_CPMDMA3LLCLK(0),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXREM_CPMDMA3LLCLK_posedge_posedge(0),
	SetupLow => tsetup_LLDMA3RXREM_CPMDMA3LLCLK_negedge_posedge(0),
	HoldLow => thold_LLDMA3RXREM_CPMDMA3LLCLK_posedge_posedge(0),
	HoldHigh => thold_LLDMA3RXREM_CPMDMA3LLCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXREM1_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXREM1_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXREM_dly(1),
	TestSignalName => "LLDMA3RXREM(1)",
	TestDelay => tisd_LLDMA3RXREM_CPMDMA3LLCLK(1),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXREM_CPMDMA3LLCLK_posedge_posedge(1),
	SetupLow => tsetup_LLDMA3RXREM_CPMDMA3LLCLK_negedge_posedge(1),
	HoldLow => thold_LLDMA3RXREM_CPMDMA3LLCLK_posedge_posedge(1),
	HoldHigh => thold_LLDMA3RXREM_CPMDMA3LLCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXREM2_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXREM2_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXREM_dly(2),
	TestSignalName => "LLDMA3RXREM(2)",
	TestDelay => tisd_LLDMA3RXREM_CPMDMA3LLCLK(2),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXREM_CPMDMA3LLCLK_posedge_posedge(2),
	SetupLow => tsetup_LLDMA3RXREM_CPMDMA3LLCLK_negedge_posedge(2),
	HoldLow => thold_LLDMA3RXREM_CPMDMA3LLCLK_posedge_posedge(2),
	HoldHigh => thold_LLDMA3RXREM_CPMDMA3LLCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_LLDMA3RXREM3_CPMDMA3LLCLK_posedge,
	TimingData => Tmkr_LLDMA3RXREM3_CPMDMA3LLCLK_posedge,
	TestSignal => LLDMA3RXREM_dly(3),
	TestSignalName => "LLDMA3RXREM(3)",
	TestDelay => tisd_LLDMA3RXREM_CPMDMA3LLCLK(3),
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName => "CPMDMA3LLCLK",
	RefDelay => ticd_CPMDMA3LLCLK,
	SetupHigh => tsetup_LLDMA3RXREM_CPMDMA3LLCLK_posedge_posedge(3),
	SetupLow => tsetup_LLDMA3RXREM_CPMDMA3LLCLK_negedge_posedge(3),
	HoldLow => thold_LLDMA3RXREM_CPMDMA3LLCLK_posedge_posedge(3),
	HoldHigh => thold_LLDMA3RXREM_CPMDMA3LLCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA3RXSOFN_CPMDMA3LLCLK_posedge,
	TimingData     => Tmkr_LLDMA3RXSOFN_CPMDMA3LLCLK_posedge,
	TestSignal     => LLDMA3RXSOFN,
	TestSignalName => "LLDMA3RXSOFN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName  => "CPMDMA3LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA3RXSOFN_CPMDMA3LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA3RXSOFN_CPMDMA3LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA3RXSOFN_CPMDMA3LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA3RXSOFN_CPMDMA3LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA3RXSOPN_CPMDMA3LLCLK_posedge,
	TimingData     => Tmkr_LLDMA3RXSOPN_CPMDMA3LLCLK_posedge,
	TestSignal     => LLDMA3RXSOPN,
	TestSignalName => "LLDMA3RXSOPN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName  => "CPMDMA3LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA3RXSOPN_CPMDMA3LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA3RXSOPN_CPMDMA3LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA3RXSOPN_CPMDMA3LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA3RXSOPN_CPMDMA3LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA3RXSRCRDYN_CPMDMA3LLCLK_posedge,
	TimingData     => Tmkr_LLDMA3RXSRCRDYN_CPMDMA3LLCLK_posedge,
	TestSignal     => LLDMA3RXSRCRDYN,
	TestSignalName => "LLDMA3RXSRCRDYN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName  => "CPMDMA3LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA3RXSRCRDYN_CPMDMA3LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA3RXSRCRDYN_CPMDMA3LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA3RXSRCRDYN_CPMDMA3LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA3RXSRCRDYN_CPMDMA3LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_LLDMA3TXDSTRDYN_CPMDMA3LLCLK_posedge,
	TimingData     => Tmkr_LLDMA3TXDSTRDYN_CPMDMA3LLCLK_posedge,
	TestSignal     => LLDMA3TXDSTRDYN,
	TestSignalName => "LLDMA3TXDSTRDYN",
	TestDelay      => 0 ps,
	RefSignal => CPMDMA3LLCLK_dly,
	RefSignalName  => "CPMDMA3LLCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_LLDMA3TXDSTRDYN_CPMDMA3LLCLK_posedge_posedge,
	SetupLow       => tsetup_LLDMA3TXDSTRDYN_CPMDMA3LLCLK_negedge_posedge,
	HoldLow        => thold_LLDMA3TXDSTRDYN_CPMDMA3LLCLK_posedge_posedge,
	HoldHigh       => thold_LLDMA3TXDSTRDYN_CPMDMA3LLCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCMADDRACK_CPMPPCMPLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCMADDRACK_CPMPPCMPLBCLK_posedge,
	TestSignal     => PLBPPCMADDRACK,
	TestSignalName => "PLBPPCMADDRACK",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName  => "CPMPPCMPLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCMADDRACK_CPMPPCMPLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCMADDRACK_CPMPPCMPLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCMADDRACK_CPMPPCMPLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCMADDRACK_CPMPPCMPLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCMMBUSY_CPMPPCMPLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCMMBUSY_CPMPPCMPLBCLK_posedge,
	TestSignal     => PLBPPCMMBUSY,
	TestSignalName => "PLBPPCMMBUSY",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName  => "CPMPPCMPLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCMMBUSY_CPMPPCMPLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCMMBUSY_CPMPPCMPLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCMMBUSY_CPMPPCMPLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCMMBUSY_CPMPPCMPLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCMMIRQ_CPMPPCMPLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCMMIRQ_CPMPPCMPLBCLK_posedge,
	TestSignal     => PLBPPCMMIRQ,
	TestSignalName => "PLBPPCMMIRQ",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName  => "CPMPPCMPLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCMMIRQ_CPMPPCMPLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCMMIRQ_CPMPPCMPLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCMMIRQ_CPMPPCMPLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCMMIRQ_CPMPPCMPLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCMMRDERR_CPMPPCMPLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCMMRDERR_CPMPPCMPLBCLK_posedge,
	TestSignal     => PLBPPCMMRDERR,
	TestSignalName => "PLBPPCMMRDERR",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName  => "CPMPPCMPLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCMMRDERR_CPMPPCMPLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCMMRDERR_CPMPPCMPLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCMMRDERR_CPMPPCMPLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCMMRDERR_CPMPPCMPLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCMMWRERR_CPMPPCMPLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCMMWRERR_CPMPPCMPLBCLK_posedge,
	TestSignal     => PLBPPCMMWRERR,
	TestSignalName => "PLBPPCMMWRERR",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName  => "CPMPPCMPLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCMMWRERR_CPMPPCMPLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCMMWRERR_CPMPPCMPLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCMMWRERR_CPMPPCMPLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCMMWRERR_CPMPPCMPLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCMRDBTERM_CPMPPCMPLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCMRDBTERM_CPMPPCMPLBCLK_posedge,
	TestSignal     => PLBPPCMRDBTERM,
	TestSignalName => "PLBPPCMRDBTERM",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName  => "CPMPPCMPLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCMRDBTERM_CPMPPCMPLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCMRDBTERM_CPMPPCMPLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCMRDBTERM_CPMPPCMPLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCMRDBTERM_CPMPPCMPLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCMRDDACK_CPMPPCMPLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCMRDDACK_CPMPPCMPLBCLK_posedge,
	TestSignal     => PLBPPCMRDDACK,
	TestSignalName => "PLBPPCMRDDACK",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName  => "CPMPPCMPLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCMRDDACK_CPMPPCMPLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCMRDDACK_CPMPPCMPLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCMRDDACK_CPMPPCMPLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCMRDDACK_CPMPPCMPLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS0_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS0_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(0),
	TestSignalName => "PLBPPCMRDDBUS(0)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(0),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS1_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS1_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(1),
	TestSignalName => "PLBPPCMRDDBUS(1)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(1),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS2_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS2_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(2),
	TestSignalName => "PLBPPCMRDDBUS(2)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(2),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(2),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(2),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(2),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS3_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS3_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(3),
	TestSignalName => "PLBPPCMRDDBUS(3)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(3),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(3),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(3),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(3),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS4_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS4_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(4),
	TestSignalName => "PLBPPCMRDDBUS(4)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(4),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(4),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(4),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(4),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS5_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS5_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(5),
	TestSignalName => "PLBPPCMRDDBUS(5)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(5),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(5),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(5),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(5),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS6_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS6_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(6),
	TestSignalName => "PLBPPCMRDDBUS(6)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(6),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(6),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(6),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(6),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS7_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS7_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(7),
	TestSignalName => "PLBPPCMRDDBUS(7)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(7),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(7),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(7),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(7),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS8_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS8_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(8),
	TestSignalName => "PLBPPCMRDDBUS(8)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(8),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(8),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(8),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(8),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS9_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS9_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(9),
	TestSignalName => "PLBPPCMRDDBUS(9)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(9),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(9),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(9),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(9),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS10_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS10_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(10),
	TestSignalName => "PLBPPCMRDDBUS(10)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(10),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(10),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(10),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(10),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS11_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS11_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(11),
	TestSignalName => "PLBPPCMRDDBUS(11)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(11),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(11),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(11),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(11),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS12_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS12_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(12),
	TestSignalName => "PLBPPCMRDDBUS(12)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(12),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(12),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(12),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(12),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS13_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS13_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(13),
	TestSignalName => "PLBPPCMRDDBUS(13)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(13),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(13),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(13),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(13),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS14_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS14_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(14),
	TestSignalName => "PLBPPCMRDDBUS(14)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(14),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(14),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(14),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(14),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS15_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS15_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(15),
	TestSignalName => "PLBPPCMRDDBUS(15)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(15),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(15),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(15),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(15),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS16_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS16_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(16),
	TestSignalName => "PLBPPCMRDDBUS(16)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(16),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(16),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(16),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(16),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(16),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS17_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS17_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(17),
	TestSignalName => "PLBPPCMRDDBUS(17)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(17),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(17),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(17),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(17),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(17),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS18_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS18_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(18),
	TestSignalName => "PLBPPCMRDDBUS(18)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(18),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(18),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(18),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(18),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(18),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS19_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS19_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(19),
	TestSignalName => "PLBPPCMRDDBUS(19)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(19),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(19),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(19),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(19),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(19),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS20_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS20_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(20),
	TestSignalName => "PLBPPCMRDDBUS(20)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(20),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(20),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(20),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(20),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(20),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS21_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS21_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(21),
	TestSignalName => "PLBPPCMRDDBUS(21)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(21),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(21),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(21),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(21),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(21),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS22_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS22_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(22),
	TestSignalName => "PLBPPCMRDDBUS(22)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(22),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(22),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(22),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(22),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(22),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS23_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS23_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(23),
	TestSignalName => "PLBPPCMRDDBUS(23)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(23),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(23),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(23),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(23),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(23),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS24_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS24_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(24),
	TestSignalName => "PLBPPCMRDDBUS(24)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(24),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(24),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(24),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(24),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(24),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS25_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS25_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(25),
	TestSignalName => "PLBPPCMRDDBUS(25)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(25),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(25),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(25),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(25),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(25),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS26_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS26_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(26),
	TestSignalName => "PLBPPCMRDDBUS(26)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(26),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(26),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(26),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(26),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(26),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS27_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS27_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(27),
	TestSignalName => "PLBPPCMRDDBUS(27)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(27),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(27),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(27),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(27),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(27),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS28_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS28_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(28),
	TestSignalName => "PLBPPCMRDDBUS(28)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(28),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(28),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(28),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(28),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS29_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS29_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(29),
	TestSignalName => "PLBPPCMRDDBUS(29)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(29),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(29),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(29),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(29),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS30_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS30_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(30),
	TestSignalName => "PLBPPCMRDDBUS(30)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(30),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(30),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(30),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(30),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS31_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS31_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(31),
	TestSignalName => "PLBPPCMRDDBUS(31)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(31),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(31),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(31),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(31),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS32_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS32_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(32),
	TestSignalName => "PLBPPCMRDDBUS(32)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(32),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(32),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(32),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(32),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(32),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS33_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS33_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(33),
	TestSignalName => "PLBPPCMRDDBUS(33)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(33),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(33),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(33),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(33),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(33),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS34_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS34_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(34),
	TestSignalName => "PLBPPCMRDDBUS(34)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(34),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(34),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(34),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(34),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(34),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS35_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS35_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(35),
	TestSignalName => "PLBPPCMRDDBUS(35)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(35),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(35),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(35),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(35),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(35),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS36_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS36_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(36),
	TestSignalName => "PLBPPCMRDDBUS(36)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(36),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(36),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(36),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(36),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(36),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS37_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS37_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(37),
	TestSignalName => "PLBPPCMRDDBUS(37)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(37),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(37),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(37),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(37),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(37),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS38_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS38_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(38),
	TestSignalName => "PLBPPCMRDDBUS(38)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(38),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(38),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(38),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(38),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(38),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS39_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS39_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(39),
	TestSignalName => "PLBPPCMRDDBUS(39)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(39),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(39),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(39),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(39),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(39),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS40_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS40_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(40),
	TestSignalName => "PLBPPCMRDDBUS(40)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(40),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(40),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(40),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(40),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(40),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS41_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS41_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(41),
	TestSignalName => "PLBPPCMRDDBUS(41)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(41),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(41),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(41),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(41),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(41),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS42_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS42_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(42),
	TestSignalName => "PLBPPCMRDDBUS(42)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(42),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(42),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(42),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(42),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(42),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS43_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS43_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(43),
	TestSignalName => "PLBPPCMRDDBUS(43)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(43),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(43),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(43),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(43),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(43),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS44_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS44_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(44),
	TestSignalName => "PLBPPCMRDDBUS(44)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(44),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(44),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(44),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(44),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(44),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS45_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS45_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(45),
	TestSignalName => "PLBPPCMRDDBUS(45)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(45),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(45),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(45),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(45),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(45),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS46_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS46_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(46),
	TestSignalName => "PLBPPCMRDDBUS(46)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(46),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(46),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(46),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(46),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(46),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS47_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS47_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(47),
	TestSignalName => "PLBPPCMRDDBUS(47)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(47),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(47),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(47),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(47),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(47),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS48_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS48_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(48),
	TestSignalName => "PLBPPCMRDDBUS(48)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(48),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(48),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(48),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(48),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(48),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS49_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS49_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(49),
	TestSignalName => "PLBPPCMRDDBUS(49)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(49),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(49),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(49),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(49),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(49),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS50_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS50_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(50),
	TestSignalName => "PLBPPCMRDDBUS(50)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(50),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(50),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(50),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(50),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(50),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS51_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS51_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(51),
	TestSignalName => "PLBPPCMRDDBUS(51)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(51),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(51),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(51),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(51),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(51),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS52_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS52_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(52),
	TestSignalName => "PLBPPCMRDDBUS(52)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(52),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(52),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(52),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(52),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(52),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS53_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS53_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(53),
	TestSignalName => "PLBPPCMRDDBUS(53)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(53),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(53),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(53),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(53),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(53),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS54_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS54_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(54),
	TestSignalName => "PLBPPCMRDDBUS(54)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(54),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(54),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(54),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(54),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(54),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS55_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS55_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(55),
	TestSignalName => "PLBPPCMRDDBUS(55)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(55),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(55),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(55),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(55),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(55),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS56_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS56_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(56),
	TestSignalName => "PLBPPCMRDDBUS(56)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(56),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(56),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(56),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(56),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(56),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS57_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS57_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(57),
	TestSignalName => "PLBPPCMRDDBUS(57)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(57),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(57),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(57),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(57),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(57),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS58_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS58_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(58),
	TestSignalName => "PLBPPCMRDDBUS(58)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(58),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(58),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(58),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(58),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(58),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS59_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS59_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(59),
	TestSignalName => "PLBPPCMRDDBUS(59)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(59),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(59),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(59),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(59),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(59),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS60_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS60_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(60),
	TestSignalName => "PLBPPCMRDDBUS(60)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(60),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(60),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(60),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(60),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(60),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS61_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS61_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(61),
	TestSignalName => "PLBPPCMRDDBUS(61)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(61),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(61),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(61),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(61),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(61),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS62_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS62_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(62),
	TestSignalName => "PLBPPCMRDDBUS(62)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(62),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(62),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(62),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(62),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(62),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS63_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS63_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(63),
	TestSignalName => "PLBPPCMRDDBUS(63)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(63),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(63),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(63),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(63),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(63),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS64_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS64_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(64),
	TestSignalName => "PLBPPCMRDDBUS(64)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(64),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(64),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(64),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(64),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(64),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS65_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS65_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(65),
	TestSignalName => "PLBPPCMRDDBUS(65)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(65),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(65),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(65),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(65),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(65),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS66_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS66_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(66),
	TestSignalName => "PLBPPCMRDDBUS(66)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(66),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(66),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(66),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(66),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(66),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS67_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS67_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(67),
	TestSignalName => "PLBPPCMRDDBUS(67)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(67),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(67),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(67),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(67),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(67),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS68_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS68_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(68),
	TestSignalName => "PLBPPCMRDDBUS(68)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(68),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(68),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(68),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(68),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(68),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS69_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS69_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(69),
	TestSignalName => "PLBPPCMRDDBUS(69)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(69),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(69),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(69),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(69),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(69),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS70_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS70_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(70),
	TestSignalName => "PLBPPCMRDDBUS(70)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(70),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(70),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(70),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(70),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(70),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS71_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS71_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(71),
	TestSignalName => "PLBPPCMRDDBUS(71)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(71),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(71),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(71),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(71),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(71),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS72_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS72_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(72),
	TestSignalName => "PLBPPCMRDDBUS(72)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(72),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(72),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(72),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(72),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(72),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS73_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS73_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(73),
	TestSignalName => "PLBPPCMRDDBUS(73)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(73),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(73),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(73),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(73),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(73),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS74_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS74_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(74),
	TestSignalName => "PLBPPCMRDDBUS(74)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(74),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(74),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(74),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(74),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(74),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS75_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS75_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(75),
	TestSignalName => "PLBPPCMRDDBUS(75)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(75),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(75),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(75),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(75),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(75),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS76_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS76_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(76),
	TestSignalName => "PLBPPCMRDDBUS(76)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(76),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(76),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(76),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(76),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(76),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS77_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS77_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(77),
	TestSignalName => "PLBPPCMRDDBUS(77)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(77),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(77),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(77),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(77),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(77),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS78_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS78_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(78),
	TestSignalName => "PLBPPCMRDDBUS(78)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(78),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(78),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(78),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(78),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(78),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS79_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS79_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(79),
	TestSignalName => "PLBPPCMRDDBUS(79)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(79),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(79),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(79),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(79),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(79),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS80_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS80_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(80),
	TestSignalName => "PLBPPCMRDDBUS(80)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(80),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(80),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(80),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(80),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(80),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS81_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS81_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(81),
	TestSignalName => "PLBPPCMRDDBUS(81)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(81),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(81),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(81),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(81),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(81),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS82_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS82_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(82),
	TestSignalName => "PLBPPCMRDDBUS(82)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(82),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(82),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(82),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(82),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(82),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS83_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS83_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(83),
	TestSignalName => "PLBPPCMRDDBUS(83)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(83),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(83),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(83),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(83),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(83),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS84_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS84_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(84),
	TestSignalName => "PLBPPCMRDDBUS(84)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(84),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(84),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(84),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(84),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(84),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS85_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS85_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(85),
	TestSignalName => "PLBPPCMRDDBUS(85)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(85),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(85),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(85),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(85),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(85),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS86_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS86_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(86),
	TestSignalName => "PLBPPCMRDDBUS(86)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(86),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(86),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(86),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(86),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(86),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS87_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS87_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(87),
	TestSignalName => "PLBPPCMRDDBUS(87)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(87),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(87),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(87),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(87),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(87),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS88_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS88_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(88),
	TestSignalName => "PLBPPCMRDDBUS(88)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(88),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(88),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(88),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(88),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(88),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS89_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS89_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(89),
	TestSignalName => "PLBPPCMRDDBUS(89)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(89),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(89),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(89),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(89),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(89),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS90_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS90_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(90),
	TestSignalName => "PLBPPCMRDDBUS(90)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(90),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(90),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(90),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(90),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(90),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS91_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS91_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(91),
	TestSignalName => "PLBPPCMRDDBUS(91)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(91),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(91),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(91),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(91),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(91),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS92_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS92_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(92),
	TestSignalName => "PLBPPCMRDDBUS(92)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(92),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(92),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(92),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(92),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(92),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS93_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS93_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(93),
	TestSignalName => "PLBPPCMRDDBUS(93)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(93),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(93),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(93),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(93),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(93),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS94_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS94_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(94),
	TestSignalName => "PLBPPCMRDDBUS(94)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(94),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(94),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(94),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(94),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(94),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS95_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS95_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(95),
	TestSignalName => "PLBPPCMRDDBUS(95)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(95),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(95),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(95),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(95),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(95),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS96_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS96_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(96),
	TestSignalName => "PLBPPCMRDDBUS(96)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(96),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(96),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(96),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(96),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(96),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS97_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS97_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(97),
	TestSignalName => "PLBPPCMRDDBUS(97)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(97),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(97),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(97),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(97),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(97),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS98_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS98_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(98),
	TestSignalName => "PLBPPCMRDDBUS(98)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(98),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(98),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(98),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(98),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(98),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS99_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS99_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(99),
	TestSignalName => "PLBPPCMRDDBUS(99)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(99),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(99),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(99),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(99),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(99),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS100_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS100_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(100),
	TestSignalName => "PLBPPCMRDDBUS(100)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(100),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(100),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(100),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(100),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(100),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS101_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS101_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(101),
	TestSignalName => "PLBPPCMRDDBUS(101)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(101),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(101),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(101),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(101),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(101),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS102_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS102_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(102),
	TestSignalName => "PLBPPCMRDDBUS(102)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(102),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(102),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(102),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(102),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(102),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS103_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS103_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(103),
	TestSignalName => "PLBPPCMRDDBUS(103)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(103),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(103),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(103),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(103),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(103),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS104_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS104_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(104),
	TestSignalName => "PLBPPCMRDDBUS(104)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(104),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(104),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(104),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(104),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(104),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS105_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS105_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(105),
	TestSignalName => "PLBPPCMRDDBUS(105)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(105),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(105),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(105),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(105),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(105),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS106_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS106_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(106),
	TestSignalName => "PLBPPCMRDDBUS(106)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(106),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(106),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(106),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(106),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(106),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS107_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS107_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(107),
	TestSignalName => "PLBPPCMRDDBUS(107)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(107),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(107),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(107),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(107),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(107),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS108_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS108_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(108),
	TestSignalName => "PLBPPCMRDDBUS(108)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(108),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(108),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(108),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(108),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(108),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS109_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS109_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(109),
	TestSignalName => "PLBPPCMRDDBUS(109)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(109),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(109),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(109),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(109),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(109),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS110_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS110_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(110),
	TestSignalName => "PLBPPCMRDDBUS(110)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(110),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(110),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(110),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(110),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(110),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS111_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS111_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(111),
	TestSignalName => "PLBPPCMRDDBUS(111)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(111),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(111),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(111),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(111),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(111),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS112_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS112_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(112),
	TestSignalName => "PLBPPCMRDDBUS(112)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(112),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(112),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(112),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(112),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(112),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS113_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS113_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(113),
	TestSignalName => "PLBPPCMRDDBUS(113)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(113),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(113),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(113),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(113),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(113),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS114_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS114_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(114),
	TestSignalName => "PLBPPCMRDDBUS(114)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(114),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(114),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(114),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(114),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(114),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS115_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS115_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(115),
	TestSignalName => "PLBPPCMRDDBUS(115)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(115),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(115),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(115),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(115),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(115),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS116_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS116_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(116),
	TestSignalName => "PLBPPCMRDDBUS(116)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(116),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(116),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(116),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(116),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(116),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS117_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS117_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(117),
	TestSignalName => "PLBPPCMRDDBUS(117)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(117),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(117),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(117),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(117),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(117),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS118_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS118_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(118),
	TestSignalName => "PLBPPCMRDDBUS(118)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(118),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(118),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(118),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(118),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(118),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS119_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS119_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(119),
	TestSignalName => "PLBPPCMRDDBUS(119)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(119),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(119),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(119),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(119),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(119),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS120_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS120_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(120),
	TestSignalName => "PLBPPCMRDDBUS(120)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(120),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(120),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(120),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(120),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(120),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS121_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS121_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(121),
	TestSignalName => "PLBPPCMRDDBUS(121)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(121),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(121),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(121),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(121),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(121),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS122_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS122_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(122),
	TestSignalName => "PLBPPCMRDDBUS(122)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(122),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(122),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(122),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(122),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(122),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS123_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS123_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(123),
	TestSignalName => "PLBPPCMRDDBUS(123)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(123),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(123),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(123),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(123),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(123),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS124_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS124_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(124),
	TestSignalName => "PLBPPCMRDDBUS(124)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(124),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(124),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(124),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(124),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(124),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS125_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS125_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(125),
	TestSignalName => "PLBPPCMRDDBUS(125)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(125),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(125),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(125),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(125),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(125),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS126_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS126_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(126),
	TestSignalName => "PLBPPCMRDDBUS(126)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(126),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(126),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(126),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(126),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(126),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDDBUS127_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDDBUS127_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDDBUS_dly(127),
	TestSignalName => "PLBPPCMRDDBUS(127)",
	TestDelay => tisd_PLBPPCMRDDBUS_CPMPPCMPLBCLK(127),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(127),
	SetupLow => tsetup_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(127),
	HoldLow => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_posedge_posedge(127),
	HoldHigh => thold_PLBPPCMRDDBUS_CPMPPCMPLBCLK_negedge_posedge(127),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDPENDPRI0_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDPENDPRI0_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDPENDPRI_dly(0),
	TestSignalName => "PLBPPCMRDPENDPRI(0)",
	TestDelay => tisd_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK(0),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDPENDPRI1_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDPENDPRI1_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDPENDPRI_dly(1),
	TestSignalName => "PLBPPCMRDPENDPRI(1)",
	TestDelay => tisd_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK(1),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCMRDPENDPRI_CPMPPCMPLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCMRDPENDREQ_CPMPPCMPLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCMRDPENDREQ_CPMPPCMPLBCLK_posedge,
	TestSignal     => PLBPPCMRDPENDREQ,
	TestSignalName => "PLBPPCMRDPENDREQ",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName  => "CPMPPCMPLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCMRDPENDREQ_CPMPPCMPLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCMRDPENDREQ_CPMPPCMPLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCMRDPENDREQ_CPMPPCMPLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCMRDPENDREQ_CPMPPCMPLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDWDADDR0_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDWDADDR0_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDWDADDR_dly(0),
	TestSignalName => "PLBPPCMRDWDADDR(0)",
	TestDelay => tisd_PLBPPCMRDWDADDR_CPMPPCMPLBCLK(0),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDWDADDR1_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDWDADDR1_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDWDADDR_dly(1),
	TestSignalName => "PLBPPCMRDWDADDR(1)",
	TestDelay => tisd_PLBPPCMRDWDADDR_CPMPPCMPLBCLK(1),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDWDADDR2_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDWDADDR2_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDWDADDR_dly(2),
	TestSignalName => "PLBPPCMRDWDADDR(2)",
	TestDelay => tisd_PLBPPCMRDWDADDR_CPMPPCMPLBCLK(2),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_posedge_posedge(2),
	SetupLow => tsetup_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_negedge_posedge(2),
	HoldLow => thold_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_posedge_posedge(2),
	HoldHigh => thold_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMRDWDADDR3_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMRDWDADDR3_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMRDWDADDR_dly(3),
	TestSignalName => "PLBPPCMRDWDADDR(3)",
	TestDelay => tisd_PLBPPCMRDWDADDR_CPMPPCMPLBCLK(3),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_posedge_posedge(3),
	SetupLow => tsetup_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_negedge_posedge(3),
	HoldLow => thold_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_posedge_posedge(3),
	HoldHigh => thold_PLBPPCMRDWDADDR_CPMPPCMPLBCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCMREARBITRATE_CPMPPCMPLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCMREARBITRATE_CPMPPCMPLBCLK_posedge,
	TestSignal     => PLBPPCMREARBITRATE,
	TestSignalName => "PLBPPCMREARBITRATE",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName  => "CPMPPCMPLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCMREARBITRATE_CPMPPCMPLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCMREARBITRATE_CPMPPCMPLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCMREARBITRATE_CPMPPCMPLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCMREARBITRATE_CPMPPCMPLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMREQPRI0_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMREQPRI0_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMREQPRI_dly(0),
	TestSignalName => "PLBPPCMREQPRI(0)",
	TestDelay => tisd_PLBPPCMREQPRI_CPMPPCMPLBCLK(0),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMREQPRI_CPMPPCMPLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCMREQPRI_CPMPPCMPLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCMREQPRI_CPMPPCMPLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCMREQPRI_CPMPPCMPLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMREQPRI1_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMREQPRI1_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMREQPRI_dly(1),
	TestSignalName => "PLBPPCMREQPRI(1)",
	TestDelay => tisd_PLBPPCMREQPRI_CPMPPCMPLBCLK(1),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMREQPRI_CPMPPCMPLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCMREQPRI_CPMPPCMPLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCMREQPRI_CPMPPCMPLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCMREQPRI_CPMPPCMPLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMSSIZE0_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMSSIZE0_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMSSIZE_dly(0),
	TestSignalName => "PLBPPCMSSIZE(0)",
	TestDelay => tisd_PLBPPCMSSIZE_CPMPPCMPLBCLK(0),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMSSIZE_CPMPPCMPLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCMSSIZE_CPMPPCMPLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCMSSIZE_CPMPPCMPLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCMSSIZE_CPMPPCMPLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMSSIZE1_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMSSIZE1_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMSSIZE_dly(1),
	TestSignalName => "PLBPPCMSSIZE(1)",
	TestDelay => tisd_PLBPPCMSSIZE_CPMPPCMPLBCLK(1),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMSSIZE_CPMPPCMPLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCMSSIZE_CPMPPCMPLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCMSSIZE_CPMPPCMPLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCMSSIZE_CPMPPCMPLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCMTIMEOUT_CPMPPCMPLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCMTIMEOUT_CPMPPCMPLBCLK_posedge,
	TestSignal     => PLBPPCMTIMEOUT,
	TestSignalName => "PLBPPCMTIMEOUT",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName  => "CPMPPCMPLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCMTIMEOUT_CPMPPCMPLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCMTIMEOUT_CPMPPCMPLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCMTIMEOUT_CPMPPCMPLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCMTIMEOUT_CPMPPCMPLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCMWRBTERM_CPMPPCMPLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCMWRBTERM_CPMPPCMPLBCLK_posedge,
	TestSignal     => PLBPPCMWRBTERM,
	TestSignalName => "PLBPPCMWRBTERM",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName  => "CPMPPCMPLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCMWRBTERM_CPMPPCMPLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCMWRBTERM_CPMPPCMPLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCMWRBTERM_CPMPPCMPLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCMWRBTERM_CPMPPCMPLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCMWRDACK_CPMPPCMPLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCMWRDACK_CPMPPCMPLBCLK_posedge,
	TestSignal     => PLBPPCMWRDACK,
	TestSignalName => "PLBPPCMWRDACK",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName  => "CPMPPCMPLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCMWRDACK_CPMPPCMPLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCMWRDACK_CPMPPCMPLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCMWRDACK_CPMPPCMPLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCMWRDACK_CPMPPCMPLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMWRPENDPRI0_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMWRPENDPRI0_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMWRPENDPRI_dly(0),
	TestSignalName => "PLBPPCMWRPENDPRI(0)",
	TestDelay => tisd_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK(0),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCMWRPENDPRI1_CPMPPCMPLBCLK_posedge,
	TimingData => Tmkr_PLBPPCMWRPENDPRI1_CPMPPCMPLBCLK_posedge,
	TestSignal => PLBPPCMWRPENDPRI_dly(1),
	TestSignalName => "PLBPPCMWRPENDPRI(1)",
	TestDelay => tisd_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK(1),
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName => "CPMPPCMPLBCLK",
	RefDelay => ticd_CPMPPCMPLBCLK,
	SetupHigh => tsetup_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCMWRPENDPRI_CPMPPCMPLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCMWRPENDREQ_CPMPPCMPLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCMWRPENDREQ_CPMPPCMPLBCLK_posedge,
	TestSignal     => PLBPPCMWRPENDREQ,
	TestSignalName => "PLBPPCMWRPENDREQ",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCMPLBCLK_dly,
	RefSignalName  => "CPMPPCMPLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCMWRPENDREQ_CPMPPCMPLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCMWRPENDREQ_CPMPPCMPLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCMWRPENDREQ_CPMPPCMPLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCMWRPENDREQ_CPMPPCMPLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS0ABORT_CPMPPCS0PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS0ABORT_CPMPPCS0PLBCLK_posedge,
	TestSignal     => PLBPPCS0ABORT,
	TestSignalName => "PLBPPCS0ABORT",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName  => "CPMPPCS0PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS0ABORT_CPMPPCS0PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS0ABORT_CPMPPCS0PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS0ABORT_CPMPPCS0PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS0ABORT_CPMPPCS0PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS0_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS0_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(0),
	TestSignalName => "PLBPPCS0ABUS(0)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(0),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS1_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS1_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(1),
	TestSignalName => "PLBPPCS0ABUS(1)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(1),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS2_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS2_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(2),
	TestSignalName => "PLBPPCS0ABUS(2)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(2),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(2),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(2),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(2),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS3_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS3_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(3),
	TestSignalName => "PLBPPCS0ABUS(3)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(3),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(3),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(3),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(3),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS4_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS4_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(4),
	TestSignalName => "PLBPPCS0ABUS(4)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(4),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(4),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(4),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(4),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS5_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS5_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(5),
	TestSignalName => "PLBPPCS0ABUS(5)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(5),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(5),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(5),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(5),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS6_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS6_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(6),
	TestSignalName => "PLBPPCS0ABUS(6)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(6),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(6),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(6),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(6),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS7_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS7_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(7),
	TestSignalName => "PLBPPCS0ABUS(7)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(7),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(7),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(7),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(7),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS8_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS8_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(8),
	TestSignalName => "PLBPPCS0ABUS(8)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(8),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(8),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(8),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(8),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS9_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS9_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(9),
	TestSignalName => "PLBPPCS0ABUS(9)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(9),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(9),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(9),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(9),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS10_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS10_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(10),
	TestSignalName => "PLBPPCS0ABUS(10)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(10),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(10),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(10),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(10),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS11_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS11_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(11),
	TestSignalName => "PLBPPCS0ABUS(11)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(11),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(11),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(11),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(11),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS12_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS12_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(12),
	TestSignalName => "PLBPPCS0ABUS(12)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(12),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(12),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(12),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(12),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS13_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS13_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(13),
	TestSignalName => "PLBPPCS0ABUS(13)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(13),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(13),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(13),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(13),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS14_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS14_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(14),
	TestSignalName => "PLBPPCS0ABUS(14)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(14),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(14),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(14),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(14),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS15_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS15_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(15),
	TestSignalName => "PLBPPCS0ABUS(15)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(15),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(15),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(15),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(15),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS16_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS16_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(16),
	TestSignalName => "PLBPPCS0ABUS(16)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(16),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(16),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(16),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(16),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(16),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS17_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS17_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(17),
	TestSignalName => "PLBPPCS0ABUS(17)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(17),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(17),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(17),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(17),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(17),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS18_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS18_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(18),
	TestSignalName => "PLBPPCS0ABUS(18)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(18),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(18),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(18),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(18),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(18),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS19_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS19_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(19),
	TestSignalName => "PLBPPCS0ABUS(19)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(19),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(19),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(19),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(19),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(19),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS20_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS20_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(20),
	TestSignalName => "PLBPPCS0ABUS(20)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(20),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(20),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(20),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(20),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(20),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS21_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS21_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(21),
	TestSignalName => "PLBPPCS0ABUS(21)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(21),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(21),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(21),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(21),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(21),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS22_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS22_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(22),
	TestSignalName => "PLBPPCS0ABUS(22)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(22),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(22),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(22),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(22),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(22),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS23_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS23_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(23),
	TestSignalName => "PLBPPCS0ABUS(23)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(23),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(23),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(23),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(23),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(23),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS24_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS24_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(24),
	TestSignalName => "PLBPPCS0ABUS(24)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(24),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(24),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(24),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(24),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(24),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS25_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS25_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(25),
	TestSignalName => "PLBPPCS0ABUS(25)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(25),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(25),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(25),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(25),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(25),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS26_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS26_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(26),
	TestSignalName => "PLBPPCS0ABUS(26)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(26),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(26),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(26),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(26),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(26),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS27_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS27_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(27),
	TestSignalName => "PLBPPCS0ABUS(27)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(27),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(27),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(27),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(27),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(27),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS28_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS28_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(28),
	TestSignalName => "PLBPPCS0ABUS(28)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(28),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(28),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(28),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(28),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS29_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS29_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(29),
	TestSignalName => "PLBPPCS0ABUS(29)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(29),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(29),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(29),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(29),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS30_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS30_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(30),
	TestSignalName => "PLBPPCS0ABUS(30)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(30),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(30),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(30),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(30),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0ABUS31_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0ABUS31_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0ABUS_dly(31),
	TestSignalName => "PLBPPCS0ABUS(31)",
	TestDelay => tisd_PLBPPCS0ABUS_CPMPPCS0PLBCLK(31),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(31),
	SetupLow => tsetup_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(31),
	HoldLow => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_posedge_posedge(31),
	HoldHigh => thold_PLBPPCS0ABUS_CPMPPCS0PLBCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE0_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE0_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(0),
	TestSignalName => "PLBPPCS0BE(0)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(0),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE1_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE1_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(1),
	TestSignalName => "PLBPPCS0BE(1)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(1),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE2_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE2_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(2),
	TestSignalName => "PLBPPCS0BE(2)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(2),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(2),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(2),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(2),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE3_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE3_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(3),
	TestSignalName => "PLBPPCS0BE(3)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(3),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(3),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(3),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(3),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE4_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE4_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(4),
	TestSignalName => "PLBPPCS0BE(4)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(4),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(4),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(4),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(4),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE5_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE5_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(5),
	TestSignalName => "PLBPPCS0BE(5)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(5),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(5),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(5),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(5),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE6_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE6_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(6),
	TestSignalName => "PLBPPCS0BE(6)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(6),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(6),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(6),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(6),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE7_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE7_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(7),
	TestSignalName => "PLBPPCS0BE(7)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(7),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(7),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(7),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(7),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE8_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE8_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(8),
	TestSignalName => "PLBPPCS0BE(8)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(8),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(8),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(8),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(8),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE9_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE9_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(9),
	TestSignalName => "PLBPPCS0BE(9)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(9),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(9),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(9),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(9),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE10_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE10_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(10),
	TestSignalName => "PLBPPCS0BE(10)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(10),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(10),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(10),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(10),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE11_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE11_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(11),
	TestSignalName => "PLBPPCS0BE(11)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(11),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(11),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(11),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(11),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE12_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE12_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(12),
	TestSignalName => "PLBPPCS0BE(12)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(12),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(12),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(12),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(12),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE13_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE13_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(13),
	TestSignalName => "PLBPPCS0BE(13)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(13),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(13),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(13),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(13),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE14_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE14_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(14),
	TestSignalName => "PLBPPCS0BE(14)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(14),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(14),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(14),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(14),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0BE15_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0BE15_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0BE_dly(15),
	TestSignalName => "PLBPPCS0BE(15)",
	TestDelay => tisd_PLBPPCS0BE_CPMPPCS0PLBCLK(15),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(15),
	SetupLow => tsetup_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(15),
	HoldLow => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_posedge_posedge(15),
	HoldHigh => thold_PLBPPCS0BE_CPMPPCS0PLBCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS0BUSLOCK_CPMPPCS0PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS0BUSLOCK_CPMPPCS0PLBCLK_posedge,
	TestSignal     => PLBPPCS0BUSLOCK,
	TestSignalName => "PLBPPCS0BUSLOCK",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName  => "CPMPPCS0PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS0BUSLOCK_CPMPPCS0PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS0BUSLOCK_CPMPPCS0PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS0BUSLOCK_CPMPPCS0PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS0BUSLOCK_CPMPPCS0PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS0LOCKERR_CPMPPCS0PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS0LOCKERR_CPMPPCS0PLBCLK_posedge,
	TestSignal     => PLBPPCS0LOCKERR,
	TestSignalName => "PLBPPCS0LOCKERR",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName  => "CPMPPCS0PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS0LOCKERR_CPMPPCS0PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS0LOCKERR_CPMPPCS0PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS0LOCKERR_CPMPPCS0PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS0LOCKERR_CPMPPCS0PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0MASTERID0_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0MASTERID0_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0MASTERID_dly(0),
	TestSignalName => "PLBPPCS0MASTERID(0)",
	TestDelay => tisd_PLBPPCS0MASTERID_CPMPPCS0PLBCLK(0),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0MASTERID_CPMPPCS0PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS0MASTERID_CPMPPCS0PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS0MASTERID_CPMPPCS0PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS0MASTERID_CPMPPCS0PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0MASTERID1_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0MASTERID1_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0MASTERID_dly(1),
	TestSignalName => "PLBPPCS0MASTERID(1)",
	TestDelay => tisd_PLBPPCS0MASTERID_CPMPPCS0PLBCLK(1),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0MASTERID_CPMPPCS0PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS0MASTERID_CPMPPCS0PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS0MASTERID_CPMPPCS0PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS0MASTERID_CPMPPCS0PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0MSIZE0_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0MSIZE0_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0MSIZE_dly(0),
	TestSignalName => "PLBPPCS0MSIZE(0)",
	TestDelay => tisd_PLBPPCS0MSIZE_CPMPPCS0PLBCLK(0),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0MSIZE_CPMPPCS0PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS0MSIZE_CPMPPCS0PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS0MSIZE_CPMPPCS0PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS0MSIZE_CPMPPCS0PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0MSIZE1_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0MSIZE1_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0MSIZE_dly(1),
	TestSignalName => "PLBPPCS0MSIZE(1)",
	TestDelay => tisd_PLBPPCS0MSIZE_CPMPPCS0PLBCLK(1),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0MSIZE_CPMPPCS0PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS0MSIZE_CPMPPCS0PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS0MSIZE_CPMPPCS0PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS0MSIZE_CPMPPCS0PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS0PAVALID_CPMPPCS0PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS0PAVALID_CPMPPCS0PLBCLK_posedge,
	TestSignal     => PLBPPCS0PAVALID,
	TestSignalName => "PLBPPCS0PAVALID",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName  => "CPMPPCS0PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS0PAVALID_CPMPPCS0PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS0PAVALID_CPMPPCS0PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS0PAVALID_CPMPPCS0PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS0PAVALID_CPMPPCS0PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS0RDBURST_CPMPPCS0PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS0RDBURST_CPMPPCS0PLBCLK_posedge,
	TestSignal     => PLBPPCS0RDBURST,
	TestSignalName => "PLBPPCS0RDBURST",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName  => "CPMPPCS0PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS0RDBURST_CPMPPCS0PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS0RDBURST_CPMPPCS0PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS0RDBURST_CPMPPCS0PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS0RDBURST_CPMPPCS0PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0RDPENDPRI0_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0RDPENDPRI0_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0RDPENDPRI_dly(0),
	TestSignalName => "PLBPPCS0RDPENDPRI(0)",
	TestDelay => tisd_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK(0),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0RDPENDPRI1_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0RDPENDPRI1_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0RDPENDPRI_dly(1),
	TestSignalName => "PLBPPCS0RDPENDPRI(1)",
	TestDelay => tisd_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK(1),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS0RDPENDPRI_CPMPPCS0PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS0RDPENDREQ_CPMPPCS0PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS0RDPENDREQ_CPMPPCS0PLBCLK_posedge,
	TestSignal     => PLBPPCS0RDPENDREQ,
	TestSignalName => "PLBPPCS0RDPENDREQ",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName  => "CPMPPCS0PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS0RDPENDREQ_CPMPPCS0PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS0RDPENDREQ_CPMPPCS0PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS0RDPENDREQ_CPMPPCS0PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS0RDPENDREQ_CPMPPCS0PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS0RDPRIM_CPMPPCS0PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS0RDPRIM_CPMPPCS0PLBCLK_posedge,
	TestSignal     => PLBPPCS0RDPRIM,
	TestSignalName => "PLBPPCS0RDPRIM",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName  => "CPMPPCS0PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS0RDPRIM_CPMPPCS0PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS0RDPRIM_CPMPPCS0PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS0RDPRIM_CPMPPCS0PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS0RDPRIM_CPMPPCS0PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0REQPRI0_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0REQPRI0_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0REQPRI_dly(0),
	TestSignalName => "PLBPPCS0REQPRI(0)",
	TestDelay => tisd_PLBPPCS0REQPRI_CPMPPCS0PLBCLK(0),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0REQPRI_CPMPPCS0PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS0REQPRI_CPMPPCS0PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS0REQPRI_CPMPPCS0PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS0REQPRI_CPMPPCS0PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0REQPRI1_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0REQPRI1_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0REQPRI_dly(1),
	TestSignalName => "PLBPPCS0REQPRI(1)",
	TestDelay => tisd_PLBPPCS0REQPRI_CPMPPCS0PLBCLK(1),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0REQPRI_CPMPPCS0PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS0REQPRI_CPMPPCS0PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS0REQPRI_CPMPPCS0PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS0REQPRI_CPMPPCS0PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS0SAVALID_CPMPPCS0PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS0SAVALID_CPMPPCS0PLBCLK_posedge,
	TestSignal     => PLBPPCS0SAVALID,
	TestSignalName => "PLBPPCS0SAVALID",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName  => "CPMPPCS0PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS0SAVALID_CPMPPCS0PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS0SAVALID_CPMPPCS0PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS0SAVALID_CPMPPCS0PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS0SAVALID_CPMPPCS0PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0SIZE0_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0SIZE0_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0SIZE_dly(0),
	TestSignalName => "PLBPPCS0SIZE(0)",
	TestDelay => tisd_PLBPPCS0SIZE_CPMPPCS0PLBCLK(0),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0SIZE_CPMPPCS0PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS0SIZE_CPMPPCS0PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS0SIZE_CPMPPCS0PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS0SIZE_CPMPPCS0PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0SIZE1_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0SIZE1_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0SIZE_dly(1),
	TestSignalName => "PLBPPCS0SIZE(1)",
	TestDelay => tisd_PLBPPCS0SIZE_CPMPPCS0PLBCLK(1),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0SIZE_CPMPPCS0PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS0SIZE_CPMPPCS0PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS0SIZE_CPMPPCS0PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS0SIZE_CPMPPCS0PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0SIZE2_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0SIZE2_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0SIZE_dly(2),
	TestSignalName => "PLBPPCS0SIZE(2)",
	TestDelay => tisd_PLBPPCS0SIZE_CPMPPCS0PLBCLK(2),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0SIZE_CPMPPCS0PLBCLK_posedge_posedge(2),
	SetupLow => tsetup_PLBPPCS0SIZE_CPMPPCS0PLBCLK_negedge_posedge(2),
	HoldLow => thold_PLBPPCS0SIZE_CPMPPCS0PLBCLK_posedge_posedge(2),
	HoldHigh => thold_PLBPPCS0SIZE_CPMPPCS0PLBCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0SIZE3_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0SIZE3_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0SIZE_dly(3),
	TestSignalName => "PLBPPCS0SIZE(3)",
	TestDelay => tisd_PLBPPCS0SIZE_CPMPPCS0PLBCLK(3),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0SIZE_CPMPPCS0PLBCLK_posedge_posedge(3),
	SetupLow => tsetup_PLBPPCS0SIZE_CPMPPCS0PLBCLK_negedge_posedge(3),
	HoldLow => thold_PLBPPCS0SIZE_CPMPPCS0PLBCLK_posedge_posedge(3),
	HoldHigh => thold_PLBPPCS0SIZE_CPMPPCS0PLBCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE0_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE0_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(0),
	TestSignalName => "PLBPPCS0TATTRIBUTE(0)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(0),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE1_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE1_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(1),
	TestSignalName => "PLBPPCS0TATTRIBUTE(1)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(1),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE2_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE2_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(2),
	TestSignalName => "PLBPPCS0TATTRIBUTE(2)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(2),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(2),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(2),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(2),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE3_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE3_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(3),
	TestSignalName => "PLBPPCS0TATTRIBUTE(3)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(3),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(3),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(3),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(3),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE4_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE4_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(4),
	TestSignalName => "PLBPPCS0TATTRIBUTE(4)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(4),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(4),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(4),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(4),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE5_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE5_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(5),
	TestSignalName => "PLBPPCS0TATTRIBUTE(5)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(5),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(5),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(5),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(5),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE6_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE6_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(6),
	TestSignalName => "PLBPPCS0TATTRIBUTE(6)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(6),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(6),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(6),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(6),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE7_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE7_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(7),
	TestSignalName => "PLBPPCS0TATTRIBUTE(7)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(7),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(7),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(7),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(7),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE8_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE8_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(8),
	TestSignalName => "PLBPPCS0TATTRIBUTE(8)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(8),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(8),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(8),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(8),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE9_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE9_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(9),
	TestSignalName => "PLBPPCS0TATTRIBUTE(9)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(9),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(9),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(9),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(9),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE10_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE10_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(10),
	TestSignalName => "PLBPPCS0TATTRIBUTE(10)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(10),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(10),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(10),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(10),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE11_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE11_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(11),
	TestSignalName => "PLBPPCS0TATTRIBUTE(11)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(11),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(11),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(11),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(11),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE12_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE12_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(12),
	TestSignalName => "PLBPPCS0TATTRIBUTE(12)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(12),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(12),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(12),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(12),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE13_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE13_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(13),
	TestSignalName => "PLBPPCS0TATTRIBUTE(13)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(13),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(13),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(13),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(13),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE14_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE14_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(14),
	TestSignalName => "PLBPPCS0TATTRIBUTE(14)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(14),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(14),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(14),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(14),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TATTRIBUTE15_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TATTRIBUTE15_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TATTRIBUTE_dly(15),
	TestSignalName => "PLBPPCS0TATTRIBUTE(15)",
	TestDelay => tisd_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK(15),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(15),
	SetupLow => tsetup_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(15),
	HoldLow => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_posedge_posedge(15),
	HoldHigh => thold_PLBPPCS0TATTRIBUTE_CPMPPCS0PLBCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TYPE0_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TYPE0_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TYPE_dly(0),
	TestSignalName => "PLBPPCS0TYPE(0)",
	TestDelay => tisd_PLBPPCS0TYPE_CPMPPCS0PLBCLK(0),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TYPE_CPMPPCS0PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS0TYPE_CPMPPCS0PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS0TYPE_CPMPPCS0PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS0TYPE_CPMPPCS0PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TYPE1_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TYPE1_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TYPE_dly(1),
	TestSignalName => "PLBPPCS0TYPE(1)",
	TestDelay => tisd_PLBPPCS0TYPE_CPMPPCS0PLBCLK(1),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TYPE_CPMPPCS0PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS0TYPE_CPMPPCS0PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS0TYPE_CPMPPCS0PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS0TYPE_CPMPPCS0PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0TYPE2_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0TYPE2_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0TYPE_dly(2),
	TestSignalName => "PLBPPCS0TYPE(2)",
	TestDelay => tisd_PLBPPCS0TYPE_CPMPPCS0PLBCLK(2),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0TYPE_CPMPPCS0PLBCLK_posedge_posedge(2),
	SetupLow => tsetup_PLBPPCS0TYPE_CPMPPCS0PLBCLK_negedge_posedge(2),
	HoldLow => thold_PLBPPCS0TYPE_CPMPPCS0PLBCLK_posedge_posedge(2),
	HoldHigh => thold_PLBPPCS0TYPE_CPMPPCS0PLBCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0UABUS28_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0UABUS28_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0UABUS_dly(28),
	TestSignalName => "PLBPPCS0UABUS(28)",
	TestDelay => tisd_PLBPPCS0UABUS_CPMPPCS0PLBCLK(28),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0UABUS_CPMPPCS0PLBCLK_posedge_posedge(28),
	SetupLow => tsetup_PLBPPCS0UABUS_CPMPPCS0PLBCLK_negedge_posedge(28),
	HoldLow => thold_PLBPPCS0UABUS_CPMPPCS0PLBCLK_posedge_posedge(28),
	HoldHigh => thold_PLBPPCS0UABUS_CPMPPCS0PLBCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0UABUS29_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0UABUS29_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0UABUS_dly(29),
	TestSignalName => "PLBPPCS0UABUS(29)",
	TestDelay => tisd_PLBPPCS0UABUS_CPMPPCS0PLBCLK(29),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0UABUS_CPMPPCS0PLBCLK_posedge_posedge(29),
	SetupLow => tsetup_PLBPPCS0UABUS_CPMPPCS0PLBCLK_negedge_posedge(29),
	HoldLow => thold_PLBPPCS0UABUS_CPMPPCS0PLBCLK_posedge_posedge(29),
	HoldHigh => thold_PLBPPCS0UABUS_CPMPPCS0PLBCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0UABUS30_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0UABUS30_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0UABUS_dly(30),
	TestSignalName => "PLBPPCS0UABUS(30)",
	TestDelay => tisd_PLBPPCS0UABUS_CPMPPCS0PLBCLK(30),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0UABUS_CPMPPCS0PLBCLK_posedge_posedge(30),
	SetupLow => tsetup_PLBPPCS0UABUS_CPMPPCS0PLBCLK_negedge_posedge(30),
	HoldLow => thold_PLBPPCS0UABUS_CPMPPCS0PLBCLK_posedge_posedge(30),
	HoldHigh => thold_PLBPPCS0UABUS_CPMPPCS0PLBCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0UABUS31_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0UABUS31_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0UABUS_dly(31),
	TestSignalName => "PLBPPCS0UABUS(31)",
	TestDelay => tisd_PLBPPCS0UABUS_CPMPPCS0PLBCLK(31),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0UABUS_CPMPPCS0PLBCLK_posedge_posedge(31),
	SetupLow => tsetup_PLBPPCS0UABUS_CPMPPCS0PLBCLK_negedge_posedge(31),
	HoldLow => thold_PLBPPCS0UABUS_CPMPPCS0PLBCLK_posedge_posedge(31),
	HoldHigh => thold_PLBPPCS0UABUS_CPMPPCS0PLBCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS0WRBURST_CPMPPCS0PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS0WRBURST_CPMPPCS0PLBCLK_posedge,
	TestSignal     => PLBPPCS0WRBURST,
	TestSignalName => "PLBPPCS0WRBURST",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName  => "CPMPPCS0PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS0WRBURST_CPMPPCS0PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS0WRBURST_CPMPPCS0PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS0WRBURST_CPMPPCS0PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS0WRBURST_CPMPPCS0PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS0_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS0_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(0),
	TestSignalName => "PLBPPCS0WRDBUS(0)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(0),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS1_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS1_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(1),
	TestSignalName => "PLBPPCS0WRDBUS(1)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(1),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS2_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS2_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(2),
	TestSignalName => "PLBPPCS0WRDBUS(2)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(2),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(2),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(2),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(2),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS3_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS3_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(3),
	TestSignalName => "PLBPPCS0WRDBUS(3)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(3),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(3),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(3),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(3),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS4_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS4_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(4),
	TestSignalName => "PLBPPCS0WRDBUS(4)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(4),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(4),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(4),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(4),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS5_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS5_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(5),
	TestSignalName => "PLBPPCS0WRDBUS(5)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(5),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(5),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(5),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(5),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS6_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS6_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(6),
	TestSignalName => "PLBPPCS0WRDBUS(6)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(6),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(6),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(6),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(6),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS7_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS7_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(7),
	TestSignalName => "PLBPPCS0WRDBUS(7)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(7),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(7),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(7),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(7),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS8_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS8_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(8),
	TestSignalName => "PLBPPCS0WRDBUS(8)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(8),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(8),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(8),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(8),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS9_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS9_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(9),
	TestSignalName => "PLBPPCS0WRDBUS(9)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(9),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(9),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(9),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(9),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS10_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS10_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(10),
	TestSignalName => "PLBPPCS0WRDBUS(10)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(10),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(10),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(10),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(10),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS11_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS11_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(11),
	TestSignalName => "PLBPPCS0WRDBUS(11)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(11),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(11),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(11),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(11),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS12_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS12_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(12),
	TestSignalName => "PLBPPCS0WRDBUS(12)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(12),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(12),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(12),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(12),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS13_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS13_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(13),
	TestSignalName => "PLBPPCS0WRDBUS(13)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(13),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(13),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(13),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(13),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS14_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS14_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(14),
	TestSignalName => "PLBPPCS0WRDBUS(14)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(14),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(14),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(14),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(14),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS15_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS15_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(15),
	TestSignalName => "PLBPPCS0WRDBUS(15)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(15),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(15),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(15),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(15),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS16_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS16_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(16),
	TestSignalName => "PLBPPCS0WRDBUS(16)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(16),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(16),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(16),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(16),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(16),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS17_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS17_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(17),
	TestSignalName => "PLBPPCS0WRDBUS(17)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(17),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(17),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(17),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(17),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(17),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS18_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS18_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(18),
	TestSignalName => "PLBPPCS0WRDBUS(18)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(18),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(18),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(18),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(18),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(18),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS19_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS19_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(19),
	TestSignalName => "PLBPPCS0WRDBUS(19)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(19),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(19),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(19),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(19),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(19),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS20_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS20_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(20),
	TestSignalName => "PLBPPCS0WRDBUS(20)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(20),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(20),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(20),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(20),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(20),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS21_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS21_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(21),
	TestSignalName => "PLBPPCS0WRDBUS(21)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(21),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(21),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(21),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(21),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(21),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS22_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS22_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(22),
	TestSignalName => "PLBPPCS0WRDBUS(22)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(22),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(22),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(22),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(22),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(22),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS23_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS23_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(23),
	TestSignalName => "PLBPPCS0WRDBUS(23)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(23),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(23),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(23),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(23),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(23),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS24_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS24_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(24),
	TestSignalName => "PLBPPCS0WRDBUS(24)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(24),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(24),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(24),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(24),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(24),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS25_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS25_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(25),
	TestSignalName => "PLBPPCS0WRDBUS(25)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(25),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(25),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(25),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(25),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(25),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS26_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS26_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(26),
	TestSignalName => "PLBPPCS0WRDBUS(26)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(26),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(26),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(26),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(26),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(26),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS27_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS27_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(27),
	TestSignalName => "PLBPPCS0WRDBUS(27)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(27),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(27),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(27),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(27),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(27),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS28_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS28_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(28),
	TestSignalName => "PLBPPCS0WRDBUS(28)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(28),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(28),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(28),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(28),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS29_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS29_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(29),
	TestSignalName => "PLBPPCS0WRDBUS(29)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(29),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(29),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(29),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(29),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS30_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS30_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(30),
	TestSignalName => "PLBPPCS0WRDBUS(30)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(30),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(30),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(30),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(30),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS31_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS31_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(31),
	TestSignalName => "PLBPPCS0WRDBUS(31)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(31),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(31),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(31),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(31),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS32_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS32_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(32),
	TestSignalName => "PLBPPCS0WRDBUS(32)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(32),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(32),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(32),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(32),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(32),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS33_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS33_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(33),
	TestSignalName => "PLBPPCS0WRDBUS(33)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(33),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(33),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(33),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(33),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(33),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS34_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS34_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(34),
	TestSignalName => "PLBPPCS0WRDBUS(34)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(34),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(34),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(34),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(34),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(34),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS35_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS35_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(35),
	TestSignalName => "PLBPPCS0WRDBUS(35)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(35),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(35),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(35),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(35),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(35),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS36_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS36_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(36),
	TestSignalName => "PLBPPCS0WRDBUS(36)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(36),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(36),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(36),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(36),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(36),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS37_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS37_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(37),
	TestSignalName => "PLBPPCS0WRDBUS(37)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(37),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(37),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(37),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(37),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(37),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS38_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS38_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(38),
	TestSignalName => "PLBPPCS0WRDBUS(38)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(38),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(38),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(38),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(38),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(38),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS39_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS39_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(39),
	TestSignalName => "PLBPPCS0WRDBUS(39)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(39),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(39),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(39),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(39),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(39),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS40_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS40_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(40),
	TestSignalName => "PLBPPCS0WRDBUS(40)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(40),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(40),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(40),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(40),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(40),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS41_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS41_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(41),
	TestSignalName => "PLBPPCS0WRDBUS(41)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(41),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(41),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(41),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(41),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(41),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS42_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS42_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(42),
	TestSignalName => "PLBPPCS0WRDBUS(42)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(42),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(42),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(42),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(42),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(42),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS43_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS43_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(43),
	TestSignalName => "PLBPPCS0WRDBUS(43)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(43),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(43),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(43),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(43),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(43),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS44_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS44_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(44),
	TestSignalName => "PLBPPCS0WRDBUS(44)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(44),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(44),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(44),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(44),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(44),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS45_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS45_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(45),
	TestSignalName => "PLBPPCS0WRDBUS(45)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(45),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(45),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(45),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(45),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(45),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS46_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS46_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(46),
	TestSignalName => "PLBPPCS0WRDBUS(46)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(46),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(46),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(46),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(46),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(46),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS47_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS47_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(47),
	TestSignalName => "PLBPPCS0WRDBUS(47)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(47),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(47),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(47),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(47),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(47),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS48_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS48_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(48),
	TestSignalName => "PLBPPCS0WRDBUS(48)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(48),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(48),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(48),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(48),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(48),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS49_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS49_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(49),
	TestSignalName => "PLBPPCS0WRDBUS(49)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(49),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(49),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(49),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(49),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(49),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS50_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS50_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(50),
	TestSignalName => "PLBPPCS0WRDBUS(50)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(50),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(50),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(50),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(50),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(50),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS51_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS51_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(51),
	TestSignalName => "PLBPPCS0WRDBUS(51)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(51),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(51),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(51),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(51),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(51),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS52_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS52_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(52),
	TestSignalName => "PLBPPCS0WRDBUS(52)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(52),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(52),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(52),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(52),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(52),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS53_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS53_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(53),
	TestSignalName => "PLBPPCS0WRDBUS(53)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(53),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(53),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(53),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(53),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(53),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS54_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS54_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(54),
	TestSignalName => "PLBPPCS0WRDBUS(54)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(54),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(54),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(54),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(54),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(54),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS55_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS55_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(55),
	TestSignalName => "PLBPPCS0WRDBUS(55)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(55),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(55),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(55),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(55),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(55),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS56_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS56_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(56),
	TestSignalName => "PLBPPCS0WRDBUS(56)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(56),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(56),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(56),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(56),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(56),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS57_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS57_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(57),
	TestSignalName => "PLBPPCS0WRDBUS(57)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(57),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(57),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(57),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(57),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(57),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS58_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS58_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(58),
	TestSignalName => "PLBPPCS0WRDBUS(58)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(58),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(58),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(58),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(58),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(58),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS59_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS59_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(59),
	TestSignalName => "PLBPPCS0WRDBUS(59)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(59),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(59),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(59),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(59),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(59),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS60_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS60_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(60),
	TestSignalName => "PLBPPCS0WRDBUS(60)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(60),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(60),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(60),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(60),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(60),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS61_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS61_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(61),
	TestSignalName => "PLBPPCS0WRDBUS(61)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(61),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(61),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(61),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(61),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(61),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS62_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS62_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(62),
	TestSignalName => "PLBPPCS0WRDBUS(62)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(62),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(62),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(62),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(62),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(62),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS63_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS63_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(63),
	TestSignalName => "PLBPPCS0WRDBUS(63)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(63),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(63),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(63),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(63),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(63),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS64_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS64_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(64),
	TestSignalName => "PLBPPCS0WRDBUS(64)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(64),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(64),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(64),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(64),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(64),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS65_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS65_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(65),
	TestSignalName => "PLBPPCS0WRDBUS(65)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(65),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(65),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(65),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(65),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(65),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS66_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS66_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(66),
	TestSignalName => "PLBPPCS0WRDBUS(66)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(66),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(66),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(66),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(66),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(66),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS67_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS67_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(67),
	TestSignalName => "PLBPPCS0WRDBUS(67)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(67),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(67),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(67),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(67),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(67),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS68_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS68_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(68),
	TestSignalName => "PLBPPCS0WRDBUS(68)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(68),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(68),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(68),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(68),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(68),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS69_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS69_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(69),
	TestSignalName => "PLBPPCS0WRDBUS(69)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(69),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(69),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(69),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(69),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(69),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS70_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS70_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(70),
	TestSignalName => "PLBPPCS0WRDBUS(70)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(70),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(70),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(70),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(70),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(70),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS71_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS71_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(71),
	TestSignalName => "PLBPPCS0WRDBUS(71)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(71),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(71),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(71),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(71),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(71),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS72_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS72_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(72),
	TestSignalName => "PLBPPCS0WRDBUS(72)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(72),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(72),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(72),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(72),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(72),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS73_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS73_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(73),
	TestSignalName => "PLBPPCS0WRDBUS(73)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(73),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(73),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(73),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(73),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(73),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS74_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS74_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(74),
	TestSignalName => "PLBPPCS0WRDBUS(74)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(74),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(74),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(74),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(74),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(74),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS75_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS75_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(75),
	TestSignalName => "PLBPPCS0WRDBUS(75)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(75),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(75),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(75),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(75),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(75),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS76_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS76_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(76),
	TestSignalName => "PLBPPCS0WRDBUS(76)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(76),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(76),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(76),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(76),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(76),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS77_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS77_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(77),
	TestSignalName => "PLBPPCS0WRDBUS(77)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(77),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(77),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(77),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(77),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(77),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS78_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS78_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(78),
	TestSignalName => "PLBPPCS0WRDBUS(78)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(78),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(78),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(78),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(78),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(78),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS79_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS79_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(79),
	TestSignalName => "PLBPPCS0WRDBUS(79)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(79),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(79),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(79),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(79),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(79),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS80_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS80_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(80),
	TestSignalName => "PLBPPCS0WRDBUS(80)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(80),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(80),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(80),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(80),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(80),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS81_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS81_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(81),
	TestSignalName => "PLBPPCS0WRDBUS(81)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(81),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(81),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(81),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(81),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(81),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS82_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS82_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(82),
	TestSignalName => "PLBPPCS0WRDBUS(82)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(82),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(82),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(82),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(82),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(82),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS83_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS83_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(83),
	TestSignalName => "PLBPPCS0WRDBUS(83)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(83),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(83),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(83),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(83),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(83),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS84_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS84_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(84),
	TestSignalName => "PLBPPCS0WRDBUS(84)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(84),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(84),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(84),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(84),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(84),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS85_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS85_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(85),
	TestSignalName => "PLBPPCS0WRDBUS(85)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(85),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(85),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(85),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(85),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(85),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS86_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS86_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(86),
	TestSignalName => "PLBPPCS0WRDBUS(86)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(86),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(86),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(86),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(86),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(86),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS87_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS87_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(87),
	TestSignalName => "PLBPPCS0WRDBUS(87)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(87),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(87),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(87),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(87),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(87),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS88_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS88_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(88),
	TestSignalName => "PLBPPCS0WRDBUS(88)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(88),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(88),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(88),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(88),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(88),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS89_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS89_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(89),
	TestSignalName => "PLBPPCS0WRDBUS(89)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(89),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(89),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(89),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(89),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(89),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS90_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS90_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(90),
	TestSignalName => "PLBPPCS0WRDBUS(90)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(90),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(90),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(90),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(90),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(90),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS91_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS91_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(91),
	TestSignalName => "PLBPPCS0WRDBUS(91)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(91),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(91),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(91),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(91),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(91),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS92_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS92_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(92),
	TestSignalName => "PLBPPCS0WRDBUS(92)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(92),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(92),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(92),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(92),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(92),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS93_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS93_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(93),
	TestSignalName => "PLBPPCS0WRDBUS(93)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(93),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(93),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(93),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(93),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(93),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS94_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS94_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(94),
	TestSignalName => "PLBPPCS0WRDBUS(94)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(94),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(94),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(94),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(94),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(94),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS95_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS95_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(95),
	TestSignalName => "PLBPPCS0WRDBUS(95)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(95),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(95),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(95),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(95),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(95),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS96_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS96_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(96),
	TestSignalName => "PLBPPCS0WRDBUS(96)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(96),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(96),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(96),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(96),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(96),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS97_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS97_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(97),
	TestSignalName => "PLBPPCS0WRDBUS(97)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(97),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(97),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(97),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(97),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(97),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS98_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS98_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(98),
	TestSignalName => "PLBPPCS0WRDBUS(98)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(98),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(98),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(98),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(98),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(98),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS99_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS99_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(99),
	TestSignalName => "PLBPPCS0WRDBUS(99)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(99),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(99),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(99),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(99),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(99),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS100_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS100_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(100),
	TestSignalName => "PLBPPCS0WRDBUS(100)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(100),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(100),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(100),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(100),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(100),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS101_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS101_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(101),
	TestSignalName => "PLBPPCS0WRDBUS(101)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(101),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(101),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(101),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(101),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(101),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS102_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS102_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(102),
	TestSignalName => "PLBPPCS0WRDBUS(102)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(102),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(102),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(102),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(102),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(102),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS103_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS103_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(103),
	TestSignalName => "PLBPPCS0WRDBUS(103)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(103),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(103),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(103),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(103),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(103),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS104_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS104_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(104),
	TestSignalName => "PLBPPCS0WRDBUS(104)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(104),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(104),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(104),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(104),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(104),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS105_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS105_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(105),
	TestSignalName => "PLBPPCS0WRDBUS(105)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(105),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(105),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(105),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(105),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(105),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS106_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS106_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(106),
	TestSignalName => "PLBPPCS0WRDBUS(106)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(106),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(106),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(106),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(106),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(106),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS107_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS107_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(107),
	TestSignalName => "PLBPPCS0WRDBUS(107)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(107),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(107),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(107),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(107),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(107),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS108_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS108_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(108),
	TestSignalName => "PLBPPCS0WRDBUS(108)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(108),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(108),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(108),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(108),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(108),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS109_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS109_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(109),
	TestSignalName => "PLBPPCS0WRDBUS(109)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(109),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(109),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(109),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(109),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(109),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS110_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS110_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(110),
	TestSignalName => "PLBPPCS0WRDBUS(110)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(110),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(110),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(110),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(110),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(110),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS111_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS111_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(111),
	TestSignalName => "PLBPPCS0WRDBUS(111)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(111),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(111),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(111),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(111),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(111),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS112_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS112_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(112),
	TestSignalName => "PLBPPCS0WRDBUS(112)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(112),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(112),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(112),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(112),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(112),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS113_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS113_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(113),
	TestSignalName => "PLBPPCS0WRDBUS(113)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(113),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(113),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(113),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(113),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(113),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS114_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS114_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(114),
	TestSignalName => "PLBPPCS0WRDBUS(114)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(114),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(114),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(114),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(114),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(114),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS115_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS115_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(115),
	TestSignalName => "PLBPPCS0WRDBUS(115)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(115),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(115),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(115),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(115),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(115),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS116_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS116_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(116),
	TestSignalName => "PLBPPCS0WRDBUS(116)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(116),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(116),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(116),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(116),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(116),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS117_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS117_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(117),
	TestSignalName => "PLBPPCS0WRDBUS(117)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(117),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(117),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(117),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(117),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(117),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS118_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS118_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(118),
	TestSignalName => "PLBPPCS0WRDBUS(118)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(118),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(118),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(118),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(118),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(118),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS119_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS119_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(119),
	TestSignalName => "PLBPPCS0WRDBUS(119)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(119),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(119),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(119),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(119),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(119),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS120_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS120_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(120),
	TestSignalName => "PLBPPCS0WRDBUS(120)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(120),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(120),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(120),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(120),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(120),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS121_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS121_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(121),
	TestSignalName => "PLBPPCS0WRDBUS(121)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(121),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(121),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(121),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(121),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(121),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS122_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS122_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(122),
	TestSignalName => "PLBPPCS0WRDBUS(122)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(122),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(122),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(122),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(122),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(122),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS123_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS123_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(123),
	TestSignalName => "PLBPPCS0WRDBUS(123)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(123),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(123),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(123),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(123),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(123),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS124_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS124_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(124),
	TestSignalName => "PLBPPCS0WRDBUS(124)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(124),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(124),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(124),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(124),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(124),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS125_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS125_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(125),
	TestSignalName => "PLBPPCS0WRDBUS(125)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(125),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(125),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(125),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(125),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(125),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS126_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS126_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(126),
	TestSignalName => "PLBPPCS0WRDBUS(126)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(126),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(126),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(126),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(126),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(126),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRDBUS127_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRDBUS127_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRDBUS_dly(127),
	TestSignalName => "PLBPPCS0WRDBUS(127)",
	TestDelay => tisd_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK(127),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(127),
	SetupLow => tsetup_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(127),
	HoldLow => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_posedge_posedge(127),
	HoldHigh => thold_PLBPPCS0WRDBUS_CPMPPCS0PLBCLK_negedge_posedge(127),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRPENDPRI0_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRPENDPRI0_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRPENDPRI_dly(0),
	TestSignalName => "PLBPPCS0WRPENDPRI(0)",
	TestDelay => tisd_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK(0),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS0WRPENDPRI1_CPMPPCS0PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS0WRPENDPRI1_CPMPPCS0PLBCLK_posedge,
	TestSignal => PLBPPCS0WRPENDPRI_dly(1),
	TestSignalName => "PLBPPCS0WRPENDPRI(1)",
	TestDelay => tisd_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK(1),
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName => "CPMPPCS0PLBCLK",
	RefDelay => ticd_CPMPPCS0PLBCLK,
	SetupHigh => tsetup_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS0WRPENDPRI_CPMPPCS0PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS0WRPENDREQ_CPMPPCS0PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS0WRPENDREQ_CPMPPCS0PLBCLK_posedge,
	TestSignal     => PLBPPCS0WRPENDREQ,
	TestSignalName => "PLBPPCS0WRPENDREQ",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName  => "CPMPPCS0PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS0WRPENDREQ_CPMPPCS0PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS0WRPENDREQ_CPMPPCS0PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS0WRPENDREQ_CPMPPCS0PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS0WRPENDREQ_CPMPPCS0PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS0WRPRIM_CPMPPCS0PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS0WRPRIM_CPMPPCS0PLBCLK_posedge,
	TestSignal     => PLBPPCS0WRPRIM,
	TestSignalName => "PLBPPCS0WRPRIM",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS0PLBCLK_dly,
	RefSignalName  => "CPMPPCS0PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS0WRPRIM_CPMPPCS0PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS0WRPRIM_CPMPPCS0PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS0WRPRIM_CPMPPCS0PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS0WRPRIM_CPMPPCS0PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS1ABORT_CPMPPCS1PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS1ABORT_CPMPPCS1PLBCLK_posedge,
	TestSignal     => PLBPPCS1ABORT,
	TestSignalName => "PLBPPCS1ABORT",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName  => "CPMPPCS1PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS1ABORT_CPMPPCS1PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS1ABORT_CPMPPCS1PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS1ABORT_CPMPPCS1PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS1ABORT_CPMPPCS1PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS0_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS0_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(0),
	TestSignalName => "PLBPPCS1ABUS(0)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(0),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS1_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS1_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(1),
	TestSignalName => "PLBPPCS1ABUS(1)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(1),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS2_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS2_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(2),
	TestSignalName => "PLBPPCS1ABUS(2)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(2),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(2),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(2),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(2),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS3_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS3_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(3),
	TestSignalName => "PLBPPCS1ABUS(3)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(3),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(3),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(3),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(3),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS4_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS4_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(4),
	TestSignalName => "PLBPPCS1ABUS(4)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(4),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(4),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(4),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(4),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS5_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS5_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(5),
	TestSignalName => "PLBPPCS1ABUS(5)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(5),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(5),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(5),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(5),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS6_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS6_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(6),
	TestSignalName => "PLBPPCS1ABUS(6)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(6),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(6),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(6),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(6),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS7_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS7_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(7),
	TestSignalName => "PLBPPCS1ABUS(7)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(7),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(7),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(7),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(7),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS8_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS8_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(8),
	TestSignalName => "PLBPPCS1ABUS(8)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(8),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(8),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(8),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(8),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS9_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS9_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(9),
	TestSignalName => "PLBPPCS1ABUS(9)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(9),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(9),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(9),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(9),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS10_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS10_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(10),
	TestSignalName => "PLBPPCS1ABUS(10)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(10),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(10),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(10),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(10),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS11_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS11_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(11),
	TestSignalName => "PLBPPCS1ABUS(11)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(11),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(11),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(11),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(11),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS12_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS12_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(12),
	TestSignalName => "PLBPPCS1ABUS(12)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(12),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(12),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(12),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(12),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS13_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS13_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(13),
	TestSignalName => "PLBPPCS1ABUS(13)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(13),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(13),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(13),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(13),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS14_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS14_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(14),
	TestSignalName => "PLBPPCS1ABUS(14)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(14),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(14),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(14),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(14),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS15_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS15_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(15),
	TestSignalName => "PLBPPCS1ABUS(15)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(15),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(15),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(15),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(15),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS16_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS16_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(16),
	TestSignalName => "PLBPPCS1ABUS(16)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(16),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(16),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(16),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(16),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(16),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS17_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS17_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(17),
	TestSignalName => "PLBPPCS1ABUS(17)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(17),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(17),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(17),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(17),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(17),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS18_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS18_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(18),
	TestSignalName => "PLBPPCS1ABUS(18)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(18),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(18),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(18),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(18),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(18),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS19_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS19_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(19),
	TestSignalName => "PLBPPCS1ABUS(19)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(19),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(19),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(19),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(19),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(19),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS20_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS20_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(20),
	TestSignalName => "PLBPPCS1ABUS(20)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(20),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(20),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(20),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(20),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(20),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS21_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS21_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(21),
	TestSignalName => "PLBPPCS1ABUS(21)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(21),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(21),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(21),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(21),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(21),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS22_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS22_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(22),
	TestSignalName => "PLBPPCS1ABUS(22)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(22),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(22),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(22),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(22),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(22),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS23_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS23_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(23),
	TestSignalName => "PLBPPCS1ABUS(23)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(23),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(23),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(23),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(23),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(23),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS24_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS24_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(24),
	TestSignalName => "PLBPPCS1ABUS(24)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(24),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(24),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(24),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(24),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(24),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS25_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS25_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(25),
	TestSignalName => "PLBPPCS1ABUS(25)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(25),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(25),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(25),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(25),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(25),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS26_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS26_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(26),
	TestSignalName => "PLBPPCS1ABUS(26)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(26),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(26),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(26),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(26),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(26),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS27_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS27_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(27),
	TestSignalName => "PLBPPCS1ABUS(27)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(27),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(27),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(27),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(27),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(27),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS28_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS28_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(28),
	TestSignalName => "PLBPPCS1ABUS(28)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(28),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(28),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(28),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(28),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS29_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS29_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(29),
	TestSignalName => "PLBPPCS1ABUS(29)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(29),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(29),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(29),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(29),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS30_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS30_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(30),
	TestSignalName => "PLBPPCS1ABUS(30)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(30),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(30),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(30),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(30),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1ABUS31_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1ABUS31_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1ABUS_dly(31),
	TestSignalName => "PLBPPCS1ABUS(31)",
	TestDelay => tisd_PLBPPCS1ABUS_CPMPPCS1PLBCLK(31),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(31),
	SetupLow => tsetup_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(31),
	HoldLow => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_posedge_posedge(31),
	HoldHigh => thold_PLBPPCS1ABUS_CPMPPCS1PLBCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE0_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE0_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(0),
	TestSignalName => "PLBPPCS1BE(0)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(0),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE1_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE1_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(1),
	TestSignalName => "PLBPPCS1BE(1)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(1),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE2_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE2_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(2),
	TestSignalName => "PLBPPCS1BE(2)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(2),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(2),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(2),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(2),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE3_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE3_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(3),
	TestSignalName => "PLBPPCS1BE(3)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(3),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(3),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(3),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(3),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE4_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE4_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(4),
	TestSignalName => "PLBPPCS1BE(4)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(4),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(4),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(4),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(4),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE5_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE5_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(5),
	TestSignalName => "PLBPPCS1BE(5)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(5),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(5),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(5),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(5),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE6_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE6_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(6),
	TestSignalName => "PLBPPCS1BE(6)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(6),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(6),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(6),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(6),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE7_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE7_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(7),
	TestSignalName => "PLBPPCS1BE(7)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(7),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(7),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(7),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(7),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE8_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE8_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(8),
	TestSignalName => "PLBPPCS1BE(8)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(8),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(8),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(8),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(8),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE9_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE9_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(9),
	TestSignalName => "PLBPPCS1BE(9)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(9),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(9),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(9),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(9),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE10_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE10_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(10),
	TestSignalName => "PLBPPCS1BE(10)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(10),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(10),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(10),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(10),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE11_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE11_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(11),
	TestSignalName => "PLBPPCS1BE(11)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(11),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(11),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(11),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(11),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE12_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE12_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(12),
	TestSignalName => "PLBPPCS1BE(12)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(12),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(12),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(12),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(12),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE13_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE13_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(13),
	TestSignalName => "PLBPPCS1BE(13)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(13),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(13),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(13),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(13),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE14_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE14_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(14),
	TestSignalName => "PLBPPCS1BE(14)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(14),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(14),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(14),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(14),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1BE15_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1BE15_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1BE_dly(15),
	TestSignalName => "PLBPPCS1BE(15)",
	TestDelay => tisd_PLBPPCS1BE_CPMPPCS1PLBCLK(15),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(15),
	SetupLow => tsetup_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(15),
	HoldLow => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_posedge_posedge(15),
	HoldHigh => thold_PLBPPCS1BE_CPMPPCS1PLBCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS1BUSLOCK_CPMPPCS1PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS1BUSLOCK_CPMPPCS1PLBCLK_posedge,
	TestSignal     => PLBPPCS1BUSLOCK,
	TestSignalName => "PLBPPCS1BUSLOCK",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName  => "CPMPPCS1PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS1BUSLOCK_CPMPPCS1PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS1BUSLOCK_CPMPPCS1PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS1BUSLOCK_CPMPPCS1PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS1BUSLOCK_CPMPPCS1PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS1LOCKERR_CPMPPCS1PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS1LOCKERR_CPMPPCS1PLBCLK_posedge,
	TestSignal     => PLBPPCS1LOCKERR,
	TestSignalName => "PLBPPCS1LOCKERR",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName  => "CPMPPCS1PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS1LOCKERR_CPMPPCS1PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS1LOCKERR_CPMPPCS1PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS1LOCKERR_CPMPPCS1PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS1LOCKERR_CPMPPCS1PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1MASTERID0_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1MASTERID0_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1MASTERID_dly(0),
	TestSignalName => "PLBPPCS1MASTERID(0)",
	TestDelay => tisd_PLBPPCS1MASTERID_CPMPPCS1PLBCLK(0),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1MASTERID_CPMPPCS1PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS1MASTERID_CPMPPCS1PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS1MASTERID_CPMPPCS1PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS1MASTERID_CPMPPCS1PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1MASTERID1_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1MASTERID1_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1MASTERID_dly(1),
	TestSignalName => "PLBPPCS1MASTERID(1)",
	TestDelay => tisd_PLBPPCS1MASTERID_CPMPPCS1PLBCLK(1),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1MASTERID_CPMPPCS1PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS1MASTERID_CPMPPCS1PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS1MASTERID_CPMPPCS1PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS1MASTERID_CPMPPCS1PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1MSIZE0_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1MSIZE0_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1MSIZE_dly(0),
	TestSignalName => "PLBPPCS1MSIZE(0)",
	TestDelay => tisd_PLBPPCS1MSIZE_CPMPPCS1PLBCLK(0),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1MSIZE_CPMPPCS1PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS1MSIZE_CPMPPCS1PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS1MSIZE_CPMPPCS1PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS1MSIZE_CPMPPCS1PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1MSIZE1_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1MSIZE1_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1MSIZE_dly(1),
	TestSignalName => "PLBPPCS1MSIZE(1)",
	TestDelay => tisd_PLBPPCS1MSIZE_CPMPPCS1PLBCLK(1),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1MSIZE_CPMPPCS1PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS1MSIZE_CPMPPCS1PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS1MSIZE_CPMPPCS1PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS1MSIZE_CPMPPCS1PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS1PAVALID_CPMPPCS1PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS1PAVALID_CPMPPCS1PLBCLK_posedge,
	TestSignal     => PLBPPCS1PAVALID,
	TestSignalName => "PLBPPCS1PAVALID",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName  => "CPMPPCS1PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS1PAVALID_CPMPPCS1PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS1PAVALID_CPMPPCS1PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS1PAVALID_CPMPPCS1PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS1PAVALID_CPMPPCS1PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS1RDBURST_CPMPPCS1PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS1RDBURST_CPMPPCS1PLBCLK_posedge,
	TestSignal     => PLBPPCS1RDBURST,
	TestSignalName => "PLBPPCS1RDBURST",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName  => "CPMPPCS1PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS1RDBURST_CPMPPCS1PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS1RDBURST_CPMPPCS1PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS1RDBURST_CPMPPCS1PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS1RDBURST_CPMPPCS1PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1RDPENDPRI0_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1RDPENDPRI0_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1RDPENDPRI_dly(0),
	TestSignalName => "PLBPPCS1RDPENDPRI(0)",
	TestDelay => tisd_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK(0),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1RDPENDPRI1_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1RDPENDPRI1_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1RDPENDPRI_dly(1),
	TestSignalName => "PLBPPCS1RDPENDPRI(1)",
	TestDelay => tisd_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK(1),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS1RDPENDPRI_CPMPPCS1PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS1RDPENDREQ_CPMPPCS1PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS1RDPENDREQ_CPMPPCS1PLBCLK_posedge,
	TestSignal     => PLBPPCS1RDPENDREQ,
	TestSignalName => "PLBPPCS1RDPENDREQ",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName  => "CPMPPCS1PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS1RDPENDREQ_CPMPPCS1PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS1RDPENDREQ_CPMPPCS1PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS1RDPENDREQ_CPMPPCS1PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS1RDPENDREQ_CPMPPCS1PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS1RDPRIM_CPMPPCS1PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS1RDPRIM_CPMPPCS1PLBCLK_posedge,
	TestSignal     => PLBPPCS1RDPRIM,
	TestSignalName => "PLBPPCS1RDPRIM",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName  => "CPMPPCS1PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS1RDPRIM_CPMPPCS1PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS1RDPRIM_CPMPPCS1PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS1RDPRIM_CPMPPCS1PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS1RDPRIM_CPMPPCS1PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1REQPRI0_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1REQPRI0_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1REQPRI_dly(0),
	TestSignalName => "PLBPPCS1REQPRI(0)",
	TestDelay => tisd_PLBPPCS1REQPRI_CPMPPCS1PLBCLK(0),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1REQPRI_CPMPPCS1PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS1REQPRI_CPMPPCS1PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS1REQPRI_CPMPPCS1PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS1REQPRI_CPMPPCS1PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1REQPRI1_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1REQPRI1_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1REQPRI_dly(1),
	TestSignalName => "PLBPPCS1REQPRI(1)",
	TestDelay => tisd_PLBPPCS1REQPRI_CPMPPCS1PLBCLK(1),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1REQPRI_CPMPPCS1PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS1REQPRI_CPMPPCS1PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS1REQPRI_CPMPPCS1PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS1REQPRI_CPMPPCS1PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS1SAVALID_CPMPPCS1PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS1SAVALID_CPMPPCS1PLBCLK_posedge,
	TestSignal     => PLBPPCS1SAVALID,
	TestSignalName => "PLBPPCS1SAVALID",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName  => "CPMPPCS1PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS1SAVALID_CPMPPCS1PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS1SAVALID_CPMPPCS1PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS1SAVALID_CPMPPCS1PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS1SAVALID_CPMPPCS1PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1SIZE0_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1SIZE0_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1SIZE_dly(0),
	TestSignalName => "PLBPPCS1SIZE(0)",
	TestDelay => tisd_PLBPPCS1SIZE_CPMPPCS1PLBCLK(0),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1SIZE_CPMPPCS1PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS1SIZE_CPMPPCS1PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS1SIZE_CPMPPCS1PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS1SIZE_CPMPPCS1PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1SIZE1_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1SIZE1_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1SIZE_dly(1),
	TestSignalName => "PLBPPCS1SIZE(1)",
	TestDelay => tisd_PLBPPCS1SIZE_CPMPPCS1PLBCLK(1),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1SIZE_CPMPPCS1PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS1SIZE_CPMPPCS1PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS1SIZE_CPMPPCS1PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS1SIZE_CPMPPCS1PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1SIZE2_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1SIZE2_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1SIZE_dly(2),
	TestSignalName => "PLBPPCS1SIZE(2)",
	TestDelay => tisd_PLBPPCS1SIZE_CPMPPCS1PLBCLK(2),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1SIZE_CPMPPCS1PLBCLK_posedge_posedge(2),
	SetupLow => tsetup_PLBPPCS1SIZE_CPMPPCS1PLBCLK_negedge_posedge(2),
	HoldLow => thold_PLBPPCS1SIZE_CPMPPCS1PLBCLK_posedge_posedge(2),
	HoldHigh => thold_PLBPPCS1SIZE_CPMPPCS1PLBCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1SIZE3_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1SIZE3_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1SIZE_dly(3),
	TestSignalName => "PLBPPCS1SIZE(3)",
	TestDelay => tisd_PLBPPCS1SIZE_CPMPPCS1PLBCLK(3),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1SIZE_CPMPPCS1PLBCLK_posedge_posedge(3),
	SetupLow => tsetup_PLBPPCS1SIZE_CPMPPCS1PLBCLK_negedge_posedge(3),
	HoldLow => thold_PLBPPCS1SIZE_CPMPPCS1PLBCLK_posedge_posedge(3),
	HoldHigh => thold_PLBPPCS1SIZE_CPMPPCS1PLBCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE0_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE0_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(0),
	TestSignalName => "PLBPPCS1TATTRIBUTE(0)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(0),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE1_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE1_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(1),
	TestSignalName => "PLBPPCS1TATTRIBUTE(1)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(1),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE2_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE2_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(2),
	TestSignalName => "PLBPPCS1TATTRIBUTE(2)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(2),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(2),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(2),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(2),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE3_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE3_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(3),
	TestSignalName => "PLBPPCS1TATTRIBUTE(3)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(3),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(3),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(3),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(3),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE4_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE4_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(4),
	TestSignalName => "PLBPPCS1TATTRIBUTE(4)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(4),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(4),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(4),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(4),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE5_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE5_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(5),
	TestSignalName => "PLBPPCS1TATTRIBUTE(5)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(5),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(5),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(5),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(5),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE6_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE6_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(6),
	TestSignalName => "PLBPPCS1TATTRIBUTE(6)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(6),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(6),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(6),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(6),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE7_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE7_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(7),
	TestSignalName => "PLBPPCS1TATTRIBUTE(7)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(7),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(7),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(7),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(7),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE8_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE8_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(8),
	TestSignalName => "PLBPPCS1TATTRIBUTE(8)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(8),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(8),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(8),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(8),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE9_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE9_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(9),
	TestSignalName => "PLBPPCS1TATTRIBUTE(9)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(9),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(9),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(9),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(9),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE10_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE10_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(10),
	TestSignalName => "PLBPPCS1TATTRIBUTE(10)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(10),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(10),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(10),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(10),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE11_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE11_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(11),
	TestSignalName => "PLBPPCS1TATTRIBUTE(11)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(11),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(11),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(11),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(11),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE12_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE12_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(12),
	TestSignalName => "PLBPPCS1TATTRIBUTE(12)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(12),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(12),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(12),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(12),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE13_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE13_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(13),
	TestSignalName => "PLBPPCS1TATTRIBUTE(13)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(13),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(13),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(13),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(13),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE14_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE14_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(14),
	TestSignalName => "PLBPPCS1TATTRIBUTE(14)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(14),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(14),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(14),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(14),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TATTRIBUTE15_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TATTRIBUTE15_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TATTRIBUTE_dly(15),
	TestSignalName => "PLBPPCS1TATTRIBUTE(15)",
	TestDelay => tisd_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK(15),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(15),
	SetupLow => tsetup_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(15),
	HoldLow => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_posedge_posedge(15),
	HoldHigh => thold_PLBPPCS1TATTRIBUTE_CPMPPCS1PLBCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TYPE0_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TYPE0_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TYPE_dly(0),
	TestSignalName => "PLBPPCS1TYPE(0)",
	TestDelay => tisd_PLBPPCS1TYPE_CPMPPCS1PLBCLK(0),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TYPE_CPMPPCS1PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS1TYPE_CPMPPCS1PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS1TYPE_CPMPPCS1PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS1TYPE_CPMPPCS1PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TYPE1_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TYPE1_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TYPE_dly(1),
	TestSignalName => "PLBPPCS1TYPE(1)",
	TestDelay => tisd_PLBPPCS1TYPE_CPMPPCS1PLBCLK(1),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TYPE_CPMPPCS1PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS1TYPE_CPMPPCS1PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS1TYPE_CPMPPCS1PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS1TYPE_CPMPPCS1PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1TYPE2_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1TYPE2_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1TYPE_dly(2),
	TestSignalName => "PLBPPCS1TYPE(2)",
	TestDelay => tisd_PLBPPCS1TYPE_CPMPPCS1PLBCLK(2),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1TYPE_CPMPPCS1PLBCLK_posedge_posedge(2),
	SetupLow => tsetup_PLBPPCS1TYPE_CPMPPCS1PLBCLK_negedge_posedge(2),
	HoldLow => thold_PLBPPCS1TYPE_CPMPPCS1PLBCLK_posedge_posedge(2),
	HoldHigh => thold_PLBPPCS1TYPE_CPMPPCS1PLBCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1UABUS28_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1UABUS28_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1UABUS_dly(28),
	TestSignalName => "PLBPPCS1UABUS(28)",
	TestDelay => tisd_PLBPPCS1UABUS_CPMPPCS1PLBCLK(28),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1UABUS_CPMPPCS1PLBCLK_posedge_posedge(28),
	SetupLow => tsetup_PLBPPCS1UABUS_CPMPPCS1PLBCLK_negedge_posedge(28),
	HoldLow => thold_PLBPPCS1UABUS_CPMPPCS1PLBCLK_posedge_posedge(28),
	HoldHigh => thold_PLBPPCS1UABUS_CPMPPCS1PLBCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1UABUS29_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1UABUS29_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1UABUS_dly(29),
	TestSignalName => "PLBPPCS1UABUS(29)",
	TestDelay => tisd_PLBPPCS1UABUS_CPMPPCS1PLBCLK(29),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1UABUS_CPMPPCS1PLBCLK_posedge_posedge(29),
	SetupLow => tsetup_PLBPPCS1UABUS_CPMPPCS1PLBCLK_negedge_posedge(29),
	HoldLow => thold_PLBPPCS1UABUS_CPMPPCS1PLBCLK_posedge_posedge(29),
	HoldHigh => thold_PLBPPCS1UABUS_CPMPPCS1PLBCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1UABUS30_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1UABUS30_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1UABUS_dly(30),
	TestSignalName => "PLBPPCS1UABUS(30)",
	TestDelay => tisd_PLBPPCS1UABUS_CPMPPCS1PLBCLK(30),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1UABUS_CPMPPCS1PLBCLK_posedge_posedge(30),
	SetupLow => tsetup_PLBPPCS1UABUS_CPMPPCS1PLBCLK_negedge_posedge(30),
	HoldLow => thold_PLBPPCS1UABUS_CPMPPCS1PLBCLK_posedge_posedge(30),
	HoldHigh => thold_PLBPPCS1UABUS_CPMPPCS1PLBCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1UABUS31_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1UABUS31_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1UABUS_dly(31),
	TestSignalName => "PLBPPCS1UABUS(31)",
	TestDelay => tisd_PLBPPCS1UABUS_CPMPPCS1PLBCLK(31),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1UABUS_CPMPPCS1PLBCLK_posedge_posedge(31),
	SetupLow => tsetup_PLBPPCS1UABUS_CPMPPCS1PLBCLK_negedge_posedge(31),
	HoldLow => thold_PLBPPCS1UABUS_CPMPPCS1PLBCLK_posedge_posedge(31),
	HoldHigh => thold_PLBPPCS1UABUS_CPMPPCS1PLBCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS1WRBURST_CPMPPCS1PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS1WRBURST_CPMPPCS1PLBCLK_posedge,
	TestSignal     => PLBPPCS1WRBURST,
	TestSignalName => "PLBPPCS1WRBURST",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName  => "CPMPPCS1PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS1WRBURST_CPMPPCS1PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS1WRBURST_CPMPPCS1PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS1WRBURST_CPMPPCS1PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS1WRBURST_CPMPPCS1PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS0_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS0_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(0),
	TestSignalName => "PLBPPCS1WRDBUS(0)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(0),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS1_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS1_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(1),
	TestSignalName => "PLBPPCS1WRDBUS(1)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(1),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS2_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS2_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(2),
	TestSignalName => "PLBPPCS1WRDBUS(2)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(2),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(2),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(2),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(2),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS3_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS3_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(3),
	TestSignalName => "PLBPPCS1WRDBUS(3)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(3),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(3),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(3),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(3),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS4_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS4_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(4),
	TestSignalName => "PLBPPCS1WRDBUS(4)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(4),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(4),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(4),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(4),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS5_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS5_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(5),
	TestSignalName => "PLBPPCS1WRDBUS(5)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(5),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(5),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(5),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(5),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS6_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS6_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(6),
	TestSignalName => "PLBPPCS1WRDBUS(6)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(6),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(6),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(6),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(6),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS7_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS7_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(7),
	TestSignalName => "PLBPPCS1WRDBUS(7)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(7),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(7),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(7),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(7),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS8_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS8_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(8),
	TestSignalName => "PLBPPCS1WRDBUS(8)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(8),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(8),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(8),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(8),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS9_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS9_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(9),
	TestSignalName => "PLBPPCS1WRDBUS(9)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(9),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(9),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(9),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(9),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS10_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS10_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(10),
	TestSignalName => "PLBPPCS1WRDBUS(10)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(10),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(10),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(10),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(10),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS11_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS11_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(11),
	TestSignalName => "PLBPPCS1WRDBUS(11)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(11),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(11),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(11),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(11),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS12_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS12_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(12),
	TestSignalName => "PLBPPCS1WRDBUS(12)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(12),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(12),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(12),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(12),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS13_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS13_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(13),
	TestSignalName => "PLBPPCS1WRDBUS(13)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(13),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(13),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(13),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(13),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS14_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS14_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(14),
	TestSignalName => "PLBPPCS1WRDBUS(14)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(14),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(14),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(14),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(14),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS15_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS15_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(15),
	TestSignalName => "PLBPPCS1WRDBUS(15)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(15),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(15),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(15),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(15),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS16_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS16_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(16),
	TestSignalName => "PLBPPCS1WRDBUS(16)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(16),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(16),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(16),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(16),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(16),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS17_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS17_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(17),
	TestSignalName => "PLBPPCS1WRDBUS(17)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(17),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(17),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(17),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(17),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(17),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS18_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS18_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(18),
	TestSignalName => "PLBPPCS1WRDBUS(18)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(18),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(18),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(18),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(18),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(18),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS19_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS19_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(19),
	TestSignalName => "PLBPPCS1WRDBUS(19)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(19),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(19),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(19),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(19),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(19),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS20_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS20_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(20),
	TestSignalName => "PLBPPCS1WRDBUS(20)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(20),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(20),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(20),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(20),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(20),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS21_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS21_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(21),
	TestSignalName => "PLBPPCS1WRDBUS(21)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(21),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(21),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(21),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(21),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(21),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS22_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS22_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(22),
	TestSignalName => "PLBPPCS1WRDBUS(22)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(22),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(22),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(22),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(22),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(22),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS23_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS23_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(23),
	TestSignalName => "PLBPPCS1WRDBUS(23)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(23),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(23),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(23),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(23),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(23),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS24_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS24_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(24),
	TestSignalName => "PLBPPCS1WRDBUS(24)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(24),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(24),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(24),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(24),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(24),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS25_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS25_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(25),
	TestSignalName => "PLBPPCS1WRDBUS(25)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(25),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(25),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(25),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(25),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(25),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS26_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS26_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(26),
	TestSignalName => "PLBPPCS1WRDBUS(26)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(26),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(26),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(26),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(26),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(26),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS27_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS27_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(27),
	TestSignalName => "PLBPPCS1WRDBUS(27)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(27),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(27),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(27),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(27),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(27),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS28_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS28_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(28),
	TestSignalName => "PLBPPCS1WRDBUS(28)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(28),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(28),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(28),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(28),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS29_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS29_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(29),
	TestSignalName => "PLBPPCS1WRDBUS(29)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(29),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(29),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(29),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(29),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS30_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS30_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(30),
	TestSignalName => "PLBPPCS1WRDBUS(30)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(30),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(30),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(30),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(30),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS31_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS31_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(31),
	TestSignalName => "PLBPPCS1WRDBUS(31)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(31),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(31),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(31),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(31),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS32_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS32_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(32),
	TestSignalName => "PLBPPCS1WRDBUS(32)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(32),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(32),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(32),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(32),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(32),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS33_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS33_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(33),
	TestSignalName => "PLBPPCS1WRDBUS(33)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(33),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(33),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(33),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(33),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(33),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS34_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS34_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(34),
	TestSignalName => "PLBPPCS1WRDBUS(34)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(34),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(34),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(34),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(34),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(34),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS35_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS35_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(35),
	TestSignalName => "PLBPPCS1WRDBUS(35)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(35),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(35),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(35),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(35),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(35),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS36_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS36_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(36),
	TestSignalName => "PLBPPCS1WRDBUS(36)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(36),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(36),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(36),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(36),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(36),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS37_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS37_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(37),
	TestSignalName => "PLBPPCS1WRDBUS(37)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(37),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(37),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(37),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(37),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(37),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS38_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS38_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(38),
	TestSignalName => "PLBPPCS1WRDBUS(38)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(38),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(38),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(38),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(38),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(38),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS39_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS39_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(39),
	TestSignalName => "PLBPPCS1WRDBUS(39)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(39),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(39),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(39),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(39),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(39),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS40_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS40_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(40),
	TestSignalName => "PLBPPCS1WRDBUS(40)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(40),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(40),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(40),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(40),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(40),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS41_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS41_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(41),
	TestSignalName => "PLBPPCS1WRDBUS(41)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(41),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(41),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(41),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(41),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(41),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS42_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS42_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(42),
	TestSignalName => "PLBPPCS1WRDBUS(42)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(42),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(42),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(42),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(42),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(42),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS43_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS43_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(43),
	TestSignalName => "PLBPPCS1WRDBUS(43)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(43),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(43),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(43),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(43),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(43),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS44_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS44_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(44),
	TestSignalName => "PLBPPCS1WRDBUS(44)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(44),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(44),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(44),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(44),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(44),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS45_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS45_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(45),
	TestSignalName => "PLBPPCS1WRDBUS(45)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(45),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(45),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(45),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(45),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(45),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS46_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS46_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(46),
	TestSignalName => "PLBPPCS1WRDBUS(46)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(46),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(46),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(46),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(46),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(46),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS47_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS47_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(47),
	TestSignalName => "PLBPPCS1WRDBUS(47)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(47),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(47),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(47),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(47),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(47),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS48_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS48_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(48),
	TestSignalName => "PLBPPCS1WRDBUS(48)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(48),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(48),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(48),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(48),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(48),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS49_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS49_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(49),
	TestSignalName => "PLBPPCS1WRDBUS(49)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(49),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(49),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(49),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(49),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(49),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS50_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS50_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(50),
	TestSignalName => "PLBPPCS1WRDBUS(50)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(50),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(50),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(50),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(50),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(50),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS51_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS51_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(51),
	TestSignalName => "PLBPPCS1WRDBUS(51)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(51),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(51),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(51),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(51),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(51),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS52_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS52_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(52),
	TestSignalName => "PLBPPCS1WRDBUS(52)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(52),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(52),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(52),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(52),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(52),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS53_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS53_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(53),
	TestSignalName => "PLBPPCS1WRDBUS(53)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(53),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(53),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(53),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(53),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(53),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS54_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS54_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(54),
	TestSignalName => "PLBPPCS1WRDBUS(54)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(54),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(54),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(54),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(54),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(54),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS55_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS55_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(55),
	TestSignalName => "PLBPPCS1WRDBUS(55)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(55),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(55),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(55),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(55),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(55),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS56_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS56_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(56),
	TestSignalName => "PLBPPCS1WRDBUS(56)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(56),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(56),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(56),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(56),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(56),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS57_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS57_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(57),
	TestSignalName => "PLBPPCS1WRDBUS(57)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(57),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(57),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(57),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(57),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(57),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS58_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS58_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(58),
	TestSignalName => "PLBPPCS1WRDBUS(58)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(58),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(58),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(58),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(58),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(58),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS59_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS59_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(59),
	TestSignalName => "PLBPPCS1WRDBUS(59)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(59),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(59),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(59),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(59),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(59),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS60_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS60_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(60),
	TestSignalName => "PLBPPCS1WRDBUS(60)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(60),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(60),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(60),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(60),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(60),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS61_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS61_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(61),
	TestSignalName => "PLBPPCS1WRDBUS(61)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(61),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(61),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(61),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(61),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(61),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS62_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS62_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(62),
	TestSignalName => "PLBPPCS1WRDBUS(62)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(62),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(62),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(62),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(62),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(62),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS63_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS63_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(63),
	TestSignalName => "PLBPPCS1WRDBUS(63)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(63),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(63),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(63),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(63),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(63),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS64_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS64_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(64),
	TestSignalName => "PLBPPCS1WRDBUS(64)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(64),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(64),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(64),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(64),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(64),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS65_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS65_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(65),
	TestSignalName => "PLBPPCS1WRDBUS(65)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(65),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(65),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(65),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(65),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(65),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS66_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS66_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(66),
	TestSignalName => "PLBPPCS1WRDBUS(66)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(66),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(66),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(66),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(66),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(66),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS67_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS67_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(67),
	TestSignalName => "PLBPPCS1WRDBUS(67)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(67),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(67),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(67),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(67),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(67),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS68_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS68_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(68),
	TestSignalName => "PLBPPCS1WRDBUS(68)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(68),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(68),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(68),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(68),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(68),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS69_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS69_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(69),
	TestSignalName => "PLBPPCS1WRDBUS(69)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(69),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(69),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(69),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(69),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(69),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS70_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS70_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(70),
	TestSignalName => "PLBPPCS1WRDBUS(70)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(70),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(70),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(70),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(70),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(70),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS71_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS71_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(71),
	TestSignalName => "PLBPPCS1WRDBUS(71)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(71),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(71),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(71),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(71),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(71),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS72_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS72_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(72),
	TestSignalName => "PLBPPCS1WRDBUS(72)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(72),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(72),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(72),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(72),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(72),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS73_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS73_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(73),
	TestSignalName => "PLBPPCS1WRDBUS(73)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(73),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(73),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(73),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(73),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(73),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS74_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS74_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(74),
	TestSignalName => "PLBPPCS1WRDBUS(74)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(74),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(74),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(74),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(74),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(74),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS75_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS75_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(75),
	TestSignalName => "PLBPPCS1WRDBUS(75)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(75),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(75),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(75),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(75),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(75),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS76_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS76_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(76),
	TestSignalName => "PLBPPCS1WRDBUS(76)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(76),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(76),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(76),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(76),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(76),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS77_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS77_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(77),
	TestSignalName => "PLBPPCS1WRDBUS(77)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(77),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(77),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(77),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(77),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(77),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS78_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS78_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(78),
	TestSignalName => "PLBPPCS1WRDBUS(78)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(78),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(78),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(78),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(78),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(78),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS79_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS79_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(79),
	TestSignalName => "PLBPPCS1WRDBUS(79)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(79),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(79),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(79),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(79),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(79),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS80_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS80_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(80),
	TestSignalName => "PLBPPCS1WRDBUS(80)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(80),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(80),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(80),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(80),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(80),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS81_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS81_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(81),
	TestSignalName => "PLBPPCS1WRDBUS(81)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(81),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(81),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(81),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(81),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(81),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS82_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS82_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(82),
	TestSignalName => "PLBPPCS1WRDBUS(82)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(82),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(82),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(82),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(82),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(82),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS83_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS83_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(83),
	TestSignalName => "PLBPPCS1WRDBUS(83)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(83),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(83),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(83),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(83),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(83),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS84_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS84_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(84),
	TestSignalName => "PLBPPCS1WRDBUS(84)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(84),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(84),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(84),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(84),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(84),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS85_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS85_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(85),
	TestSignalName => "PLBPPCS1WRDBUS(85)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(85),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(85),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(85),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(85),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(85),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS86_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS86_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(86),
	TestSignalName => "PLBPPCS1WRDBUS(86)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(86),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(86),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(86),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(86),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(86),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS87_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS87_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(87),
	TestSignalName => "PLBPPCS1WRDBUS(87)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(87),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(87),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(87),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(87),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(87),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS88_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS88_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(88),
	TestSignalName => "PLBPPCS1WRDBUS(88)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(88),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(88),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(88),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(88),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(88),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS89_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS89_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(89),
	TestSignalName => "PLBPPCS1WRDBUS(89)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(89),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(89),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(89),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(89),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(89),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS90_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS90_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(90),
	TestSignalName => "PLBPPCS1WRDBUS(90)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(90),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(90),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(90),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(90),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(90),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS91_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS91_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(91),
	TestSignalName => "PLBPPCS1WRDBUS(91)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(91),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(91),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(91),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(91),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(91),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS92_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS92_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(92),
	TestSignalName => "PLBPPCS1WRDBUS(92)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(92),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(92),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(92),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(92),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(92),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS93_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS93_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(93),
	TestSignalName => "PLBPPCS1WRDBUS(93)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(93),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(93),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(93),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(93),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(93),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS94_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS94_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(94),
	TestSignalName => "PLBPPCS1WRDBUS(94)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(94),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(94),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(94),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(94),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(94),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS95_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS95_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(95),
	TestSignalName => "PLBPPCS1WRDBUS(95)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(95),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(95),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(95),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(95),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(95),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS96_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS96_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(96),
	TestSignalName => "PLBPPCS1WRDBUS(96)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(96),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(96),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(96),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(96),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(96),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS97_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS97_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(97),
	TestSignalName => "PLBPPCS1WRDBUS(97)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(97),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(97),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(97),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(97),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(97),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS98_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS98_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(98),
	TestSignalName => "PLBPPCS1WRDBUS(98)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(98),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(98),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(98),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(98),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(98),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS99_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS99_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(99),
	TestSignalName => "PLBPPCS1WRDBUS(99)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(99),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(99),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(99),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(99),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(99),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS100_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS100_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(100),
	TestSignalName => "PLBPPCS1WRDBUS(100)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(100),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(100),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(100),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(100),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(100),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS101_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS101_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(101),
	TestSignalName => "PLBPPCS1WRDBUS(101)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(101),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(101),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(101),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(101),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(101),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS102_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS102_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(102),
	TestSignalName => "PLBPPCS1WRDBUS(102)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(102),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(102),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(102),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(102),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(102),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS103_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS103_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(103),
	TestSignalName => "PLBPPCS1WRDBUS(103)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(103),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(103),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(103),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(103),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(103),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS104_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS104_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(104),
	TestSignalName => "PLBPPCS1WRDBUS(104)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(104),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(104),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(104),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(104),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(104),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS105_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS105_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(105),
	TestSignalName => "PLBPPCS1WRDBUS(105)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(105),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(105),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(105),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(105),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(105),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS106_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS106_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(106),
	TestSignalName => "PLBPPCS1WRDBUS(106)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(106),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(106),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(106),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(106),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(106),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS107_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS107_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(107),
	TestSignalName => "PLBPPCS1WRDBUS(107)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(107),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(107),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(107),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(107),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(107),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS108_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS108_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(108),
	TestSignalName => "PLBPPCS1WRDBUS(108)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(108),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(108),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(108),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(108),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(108),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS109_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS109_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(109),
	TestSignalName => "PLBPPCS1WRDBUS(109)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(109),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(109),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(109),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(109),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(109),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS110_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS110_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(110),
	TestSignalName => "PLBPPCS1WRDBUS(110)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(110),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(110),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(110),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(110),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(110),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS111_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS111_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(111),
	TestSignalName => "PLBPPCS1WRDBUS(111)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(111),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(111),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(111),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(111),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(111),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS112_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS112_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(112),
	TestSignalName => "PLBPPCS1WRDBUS(112)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(112),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(112),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(112),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(112),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(112),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS113_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS113_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(113),
	TestSignalName => "PLBPPCS1WRDBUS(113)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(113),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(113),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(113),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(113),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(113),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS114_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS114_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(114),
	TestSignalName => "PLBPPCS1WRDBUS(114)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(114),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(114),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(114),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(114),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(114),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS115_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS115_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(115),
	TestSignalName => "PLBPPCS1WRDBUS(115)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(115),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(115),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(115),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(115),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(115),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS116_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS116_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(116),
	TestSignalName => "PLBPPCS1WRDBUS(116)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(116),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(116),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(116),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(116),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(116),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS117_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS117_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(117),
	TestSignalName => "PLBPPCS1WRDBUS(117)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(117),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(117),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(117),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(117),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(117),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS118_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS118_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(118),
	TestSignalName => "PLBPPCS1WRDBUS(118)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(118),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(118),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(118),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(118),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(118),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS119_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS119_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(119),
	TestSignalName => "PLBPPCS1WRDBUS(119)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(119),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(119),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(119),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(119),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(119),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS120_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS120_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(120),
	TestSignalName => "PLBPPCS1WRDBUS(120)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(120),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(120),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(120),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(120),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(120),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS121_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS121_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(121),
	TestSignalName => "PLBPPCS1WRDBUS(121)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(121),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(121),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(121),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(121),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(121),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS122_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS122_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(122),
	TestSignalName => "PLBPPCS1WRDBUS(122)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(122),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(122),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(122),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(122),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(122),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS123_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS123_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(123),
	TestSignalName => "PLBPPCS1WRDBUS(123)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(123),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(123),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(123),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(123),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(123),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS124_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS124_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(124),
	TestSignalName => "PLBPPCS1WRDBUS(124)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(124),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(124),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(124),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(124),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(124),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS125_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS125_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(125),
	TestSignalName => "PLBPPCS1WRDBUS(125)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(125),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(125),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(125),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(125),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(125),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS126_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS126_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(126),
	TestSignalName => "PLBPPCS1WRDBUS(126)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(126),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(126),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(126),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(126),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(126),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRDBUS127_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRDBUS127_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRDBUS_dly(127),
	TestSignalName => "PLBPPCS1WRDBUS(127)",
	TestDelay => tisd_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK(127),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(127),
	SetupLow => tsetup_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(127),
	HoldLow => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_posedge_posedge(127),
	HoldHigh => thold_PLBPPCS1WRDBUS_CPMPPCS1PLBCLK_negedge_posedge(127),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRPENDPRI0_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRPENDPRI0_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRPENDPRI_dly(0),
	TestSignalName => "PLBPPCS1WRPENDPRI(0)",
	TestDelay => tisd_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK(0),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK_posedge_posedge(0),
	SetupLow => tsetup_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK_negedge_posedge(0),
	HoldLow => thold_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK_posedge_posedge(0),
	HoldHigh => thold_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_PLBPPCS1WRPENDPRI1_CPMPPCS1PLBCLK_posedge,
	TimingData => Tmkr_PLBPPCS1WRPENDPRI1_CPMPPCS1PLBCLK_posedge,
	TestSignal => PLBPPCS1WRPENDPRI_dly(1),
	TestSignalName => "PLBPPCS1WRPENDPRI(1)",
	TestDelay => tisd_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK(1),
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName => "CPMPPCS1PLBCLK",
	RefDelay => ticd_CPMPPCS1PLBCLK,
	SetupHigh => tsetup_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK_posedge_posedge(1),
	SetupLow => tsetup_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK_negedge_posedge(1),
	HoldLow => thold_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK_posedge_posedge(1),
	HoldHigh => thold_PLBPPCS1WRPENDPRI_CPMPPCS1PLBCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS1WRPENDREQ_CPMPPCS1PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS1WRPENDREQ_CPMPPCS1PLBCLK_posedge,
	TestSignal     => PLBPPCS1WRPENDREQ,
	TestSignalName => "PLBPPCS1WRPENDREQ",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName  => "CPMPPCS1PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS1WRPENDREQ_CPMPPCS1PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS1WRPENDREQ_CPMPPCS1PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS1WRPENDREQ_CPMPPCS1PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS1WRPENDREQ_CPMPPCS1PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_PLBPPCS1WRPRIM_CPMPPCS1PLBCLK_posedge,
	TimingData     => Tmkr_PLBPPCS1WRPRIM_CPMPPCS1PLBCLK_posedge,
	TestSignal     => PLBPPCS1WRPRIM,
	TestSignalName => "PLBPPCS1WRPRIM",
	TestDelay      => 0 ps,
	RefSignal => CPMPPCS1PLBCLK_dly,
	RefSignalName  => "CPMPPCS1PLBCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_PLBPPCS1WRPRIM_CPMPPCS1PLBCLK_posedge_posedge,
	SetupLow       => tsetup_PLBPPCS1WRPRIM_CPMPPCS1PLBCLK_negedge_posedge,
	HoldLow        => thold_PLBPPCS1WRPRIM_CPMPPCS1PLBCLK_posedge_posedge,
	HoldHigh       => thold_PLBPPCS1WRPRIM_CPMPPCS1PLBCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_CPMC440CORECLOCKINACTIVE_JTGC440TCK_posedge,
	TimingData     => Tmkr_CPMC440CORECLOCKINACTIVE_JTGC440TCK_posedge,
	TestSignal     => CPMC440CORECLOCKINACTIVE,
	TestSignalName => "CPMC440CORECLOCKINACTIVE",
	TestDelay      => 0 ps,
	RefSignal => JTGC440TCK_dly,
	RefSignalName  => "JTGC440TCK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_CPMC440CORECLOCKINACTIVE_JTGC440TCK_posedge_posedge,
	SetupLow       => tsetup_CPMC440CORECLOCKINACTIVE_JTGC440TCK_negedge_posedge,
	HoldLow        => thold_CPMC440CORECLOCKINACTIVE_JTGC440TCK_posedge_posedge,
	HoldHigh       => thold_CPMC440CORECLOCKINACTIVE_JTGC440TCK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_DBGC440DEBUGHALT_CPMC440CLK_posedge,
	TimingData     => Tmkr_DBGC440DEBUGHALT_CPMC440CLK_posedge,
	TestSignal     => DBGC440DEBUGHALT,
	TestSignalName => "DBGC440DEBUGHALT",
	TestDelay      => 0 ps,
	RefSignal => CPMC440CLK_dly,
	RefSignalName  => "CPMC440CLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_DBGC440DEBUGHALT_CPMC440CLK_posedge_posedge,
	SetupLow       => tsetup_DBGC440DEBUGHALT_CPMC440CLK_negedge_posedge,
	HoldLow        => thold_DBGC440DEBUGHALT_CPMC440CLK_posedge_posedge,
	HoldHigh       => thold_DBGC440DEBUGHALT_CPMC440CLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DBGC440SYSTEMSTATUS0_JTGC440TCK_posedge,
	TimingData => Tmkr_DBGC440SYSTEMSTATUS0_JTGC440TCK_posedge,
	TestSignal => DBGC440SYSTEMSTATUS_dly(0),
	TestSignalName => "DBGC440SYSTEMSTATUS(0)",
	TestDelay => tisd_DBGC440SYSTEMSTATUS_JTGC440TCK(0),
	RefSignal => JTGC440TCK_dly,
	RefSignalName => "JTGC440TCK",
	RefDelay => ticd_JTGC440TCK,
	SetupHigh => tsetup_DBGC440SYSTEMSTATUS_JTGC440TCK_posedge_posedge(0),
	SetupLow => tsetup_DBGC440SYSTEMSTATUS_JTGC440TCK_negedge_posedge(0),
	HoldLow => thold_DBGC440SYSTEMSTATUS_JTGC440TCK_posedge_posedge(0),
	HoldHigh => thold_DBGC440SYSTEMSTATUS_JTGC440TCK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DBGC440SYSTEMSTATUS1_JTGC440TCK_posedge,
	TimingData => Tmkr_DBGC440SYSTEMSTATUS1_JTGC440TCK_posedge,
	TestSignal => DBGC440SYSTEMSTATUS_dly(1),
	TestSignalName => "DBGC440SYSTEMSTATUS(1)",
	TestDelay => tisd_DBGC440SYSTEMSTATUS_JTGC440TCK(1),
	RefSignal => JTGC440TCK_dly,
	RefSignalName => "JTGC440TCK",
	RefDelay => ticd_JTGC440TCK,
	SetupHigh => tsetup_DBGC440SYSTEMSTATUS_JTGC440TCK_posedge_posedge(1),
	SetupLow => tsetup_DBGC440SYSTEMSTATUS_JTGC440TCK_negedge_posedge(1),
	HoldLow => thold_DBGC440SYSTEMSTATUS_JTGC440TCK_posedge_posedge(1),
	HoldHigh => thold_DBGC440SYSTEMSTATUS_JTGC440TCK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DBGC440SYSTEMSTATUS2_JTGC440TCK_posedge,
	TimingData => Tmkr_DBGC440SYSTEMSTATUS2_JTGC440TCK_posedge,
	TestSignal => DBGC440SYSTEMSTATUS_dly(2),
	TestSignalName => "DBGC440SYSTEMSTATUS(2)",
	TestDelay => tisd_DBGC440SYSTEMSTATUS_JTGC440TCK(2),
	RefSignal => JTGC440TCK_dly,
	RefSignalName => "JTGC440TCK",
	RefDelay => ticd_JTGC440TCK,
	SetupHigh => tsetup_DBGC440SYSTEMSTATUS_JTGC440TCK_posedge_posedge(2),
	SetupLow => tsetup_DBGC440SYSTEMSTATUS_JTGC440TCK_negedge_posedge(2),
	HoldLow => thold_DBGC440SYSTEMSTATUS_JTGC440TCK_posedge_posedge(2),
	HoldHigh => thold_DBGC440SYSTEMSTATUS_JTGC440TCK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DBGC440SYSTEMSTATUS3_JTGC440TCK_posedge,
	TimingData => Tmkr_DBGC440SYSTEMSTATUS3_JTGC440TCK_posedge,
	TestSignal => DBGC440SYSTEMSTATUS_dly(3),
	TestSignalName => "DBGC440SYSTEMSTATUS(3)",
	TestDelay => tisd_DBGC440SYSTEMSTATUS_JTGC440TCK(3),
	RefSignal => JTGC440TCK_dly,
	RefSignalName => "JTGC440TCK",
	RefDelay => ticd_JTGC440TCK,
	SetupHigh => tsetup_DBGC440SYSTEMSTATUS_JTGC440TCK_posedge_posedge(3),
	SetupLow => tsetup_DBGC440SYSTEMSTATUS_JTGC440TCK_negedge_posedge(3),
	HoldLow => thold_DBGC440SYSTEMSTATUS_JTGC440TCK_posedge_posedge(3),
	HoldHigh => thold_DBGC440SYSTEMSTATUS_JTGC440TCK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DBGC440SYSTEMSTATUS4_JTGC440TCK_posedge,
	TimingData => Tmkr_DBGC440SYSTEMSTATUS4_JTGC440TCK_posedge,
	TestSignal => DBGC440SYSTEMSTATUS_dly(4),
	TestSignalName => "DBGC440SYSTEMSTATUS(4)",
	TestDelay => tisd_DBGC440SYSTEMSTATUS_JTGC440TCK(4),
	RefSignal => JTGC440TCK_dly,
	RefSignalName => "JTGC440TCK",
	RefDelay => ticd_JTGC440TCK,
	SetupHigh => tsetup_DBGC440SYSTEMSTATUS_JTGC440TCK_posedge_posedge(4),
	SetupLow => tsetup_DBGC440SYSTEMSTATUS_JTGC440TCK_negedge_posedge(4),
	HoldLow => thold_DBGC440SYSTEMSTATUS_JTGC440TCK_posedge_posedge(4),
	HoldHigh => thold_DBGC440SYSTEMSTATUS_JTGC440TCK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_DBGC440UNCONDDEBUGEVENT_CPMC440CLK_posedge,
	TimingData     => Tmkr_DBGC440UNCONDDEBUGEVENT_CPMC440CLK_posedge,
	TestSignal     => DBGC440UNCONDDEBUGEVENT,
	TestSignalName => "DBGC440UNCONDDEBUGEVENT",
	TestDelay      => 0 ps,
	RefSignal => CPMC440CLK_dly,
	RefSignalName  => "CPMC440CLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_DBGC440UNCONDDEBUGEVENT_CPMC440CLK_posedge_posedge,
	SetupLow       => tsetup_DBGC440UNCONDDEBUGEVENT_CPMC440CLK_negedge_posedge,
	HoldLow        => thold_DBGC440UNCONDDEBUGEVENT_CPMC440CLK_posedge_posedge,
	HoldHigh       => thold_DBGC440UNCONDDEBUGEVENT_CPMC440CLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSABUS0_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSABUS0_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSABUS_dly(0),
	TestSignalName => "DCRPPCDSABUS(0)",
	TestDelay => tisd_DCRPPCDSABUS_CPMDCRCLK(0),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(0),
	SetupLow => tsetup_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(0),
	HoldLow => thold_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(0),
	HoldHigh => thold_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSABUS1_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSABUS1_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSABUS_dly(1),
	TestSignalName => "DCRPPCDSABUS(1)",
	TestDelay => tisd_DCRPPCDSABUS_CPMDCRCLK(1),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(1),
	SetupLow => tsetup_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(1),
	HoldLow => thold_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(1),
	HoldHigh => thold_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSABUS2_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSABUS2_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSABUS_dly(2),
	TestSignalName => "DCRPPCDSABUS(2)",
	TestDelay => tisd_DCRPPCDSABUS_CPMDCRCLK(2),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(2),
	SetupLow => tsetup_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(2),
	HoldLow => thold_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(2),
	HoldHigh => thold_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSABUS3_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSABUS3_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSABUS_dly(3),
	TestSignalName => "DCRPPCDSABUS(3)",
	TestDelay => tisd_DCRPPCDSABUS_CPMDCRCLK(3),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(3),
	SetupLow => tsetup_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(3),
	HoldLow => thold_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(3),
	HoldHigh => thold_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSABUS4_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSABUS4_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSABUS_dly(4),
	TestSignalName => "DCRPPCDSABUS(4)",
	TestDelay => tisd_DCRPPCDSABUS_CPMDCRCLK(4),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(4),
	SetupLow => tsetup_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(4),
	HoldLow => thold_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(4),
	HoldHigh => thold_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSABUS5_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSABUS5_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSABUS_dly(5),
	TestSignalName => "DCRPPCDSABUS(5)",
	TestDelay => tisd_DCRPPCDSABUS_CPMDCRCLK(5),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(5),
	SetupLow => tsetup_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(5),
	HoldLow => thold_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(5),
	HoldHigh => thold_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSABUS6_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSABUS6_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSABUS_dly(6),
	TestSignalName => "DCRPPCDSABUS(6)",
	TestDelay => tisd_DCRPPCDSABUS_CPMDCRCLK(6),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(6),
	SetupLow => tsetup_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(6),
	HoldLow => thold_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(6),
	HoldHigh => thold_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSABUS7_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSABUS7_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSABUS_dly(7),
	TestSignalName => "DCRPPCDSABUS(7)",
	TestDelay => tisd_DCRPPCDSABUS_CPMDCRCLK(7),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(7),
	SetupLow => tsetup_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(7),
	HoldLow => thold_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(7),
	HoldHigh => thold_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSABUS8_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSABUS8_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSABUS_dly(8),
	TestSignalName => "DCRPPCDSABUS(8)",
	TestDelay => tisd_DCRPPCDSABUS_CPMDCRCLK(8),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(8),
	SetupLow => tsetup_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(8),
	HoldLow => thold_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(8),
	HoldHigh => thold_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSABUS9_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSABUS9_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSABUS_dly(9),
	TestSignalName => "DCRPPCDSABUS(9)",
	TestDelay => tisd_DCRPPCDSABUS_CPMDCRCLK(9),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(9),
	SetupLow => tsetup_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(9),
	HoldLow => thold_DCRPPCDSABUS_CPMDCRCLK_posedge_posedge(9),
	HoldHigh => thold_DCRPPCDSABUS_CPMDCRCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT0_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT0_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(0),
	TestSignalName => "DCRPPCDSDBUSOUT(0)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(0),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(0),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(0),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(0),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT1_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT1_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(1),
	TestSignalName => "DCRPPCDSDBUSOUT(1)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(1),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(1),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(1),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(1),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT2_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT2_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(2),
	TestSignalName => "DCRPPCDSDBUSOUT(2)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(2),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(2),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(2),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(2),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT3_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT3_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(3),
	TestSignalName => "DCRPPCDSDBUSOUT(3)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(3),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(3),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(3),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(3),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT4_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT4_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(4),
	TestSignalName => "DCRPPCDSDBUSOUT(4)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(4),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(4),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(4),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(4),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT5_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT5_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(5),
	TestSignalName => "DCRPPCDSDBUSOUT(5)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(5),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(5),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(5),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(5),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT6_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT6_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(6),
	TestSignalName => "DCRPPCDSDBUSOUT(6)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(6),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(6),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(6),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(6),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT7_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT7_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(7),
	TestSignalName => "DCRPPCDSDBUSOUT(7)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(7),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(7),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(7),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(7),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT8_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT8_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(8),
	TestSignalName => "DCRPPCDSDBUSOUT(8)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(8),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(8),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(8),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(8),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT9_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT9_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(9),
	TestSignalName => "DCRPPCDSDBUSOUT(9)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(9),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(9),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(9),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(9),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT10_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT10_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(10),
	TestSignalName => "DCRPPCDSDBUSOUT(10)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(10),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(10),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(10),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(10),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT11_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT11_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(11),
	TestSignalName => "DCRPPCDSDBUSOUT(11)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(11),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(11),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(11),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(11),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT12_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT12_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(12),
	TestSignalName => "DCRPPCDSDBUSOUT(12)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(12),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(12),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(12),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(12),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT13_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT13_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(13),
	TestSignalName => "DCRPPCDSDBUSOUT(13)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(13),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(13),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(13),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(13),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT14_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT14_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(14),
	TestSignalName => "DCRPPCDSDBUSOUT(14)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(14),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(14),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(14),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(14),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT15_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT15_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(15),
	TestSignalName => "DCRPPCDSDBUSOUT(15)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(15),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(15),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(15),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(15),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT16_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT16_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(16),
	TestSignalName => "DCRPPCDSDBUSOUT(16)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(16),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(16),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(16),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(16),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(16),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT17_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT17_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(17),
	TestSignalName => "DCRPPCDSDBUSOUT(17)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(17),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(17),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(17),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(17),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(17),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT18_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT18_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(18),
	TestSignalName => "DCRPPCDSDBUSOUT(18)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(18),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(18),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(18),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(18),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(18),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT19_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT19_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(19),
	TestSignalName => "DCRPPCDSDBUSOUT(19)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(19),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(19),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(19),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(19),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(19),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT20_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT20_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(20),
	TestSignalName => "DCRPPCDSDBUSOUT(20)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(20),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(20),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(20),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(20),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(20),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT21_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT21_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(21),
	TestSignalName => "DCRPPCDSDBUSOUT(21)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(21),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(21),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(21),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(21),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(21),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT22_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT22_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(22),
	TestSignalName => "DCRPPCDSDBUSOUT(22)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(22),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(22),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(22),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(22),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(22),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT23_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT23_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(23),
	TestSignalName => "DCRPPCDSDBUSOUT(23)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(23),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(23),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(23),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(23),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(23),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT24_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT24_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(24),
	TestSignalName => "DCRPPCDSDBUSOUT(24)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(24),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(24),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(24),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(24),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(24),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT25_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT25_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(25),
	TestSignalName => "DCRPPCDSDBUSOUT(25)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(25),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(25),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(25),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(25),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(25),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT26_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT26_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(26),
	TestSignalName => "DCRPPCDSDBUSOUT(26)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(26),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(26),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(26),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(26),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(26),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT27_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT27_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(27),
	TestSignalName => "DCRPPCDSDBUSOUT(27)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(27),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(27),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(27),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(27),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(27),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT28_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT28_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(28),
	TestSignalName => "DCRPPCDSDBUSOUT(28)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(28),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(28),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(28),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(28),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT29_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT29_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(29),
	TestSignalName => "DCRPPCDSDBUSOUT(29)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(29),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(29),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(29),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(29),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT30_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT30_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(30),
	TestSignalName => "DCRPPCDSDBUSOUT(30)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(30),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(30),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(30),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(30),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_DCRPPCDSDBUSOUT31_CPMDCRCLK_posedge,
	TimingData => Tmkr_DCRPPCDSDBUSOUT31_CPMDCRCLK_posedge,
	TestSignal => DCRPPCDSDBUSOUT_dly(31),
	TestSignalName => "DCRPPCDSDBUSOUT(31)",
	TestDelay => tisd_DCRPPCDSDBUSOUT_CPMDCRCLK(31),
	RefSignal => CPMDCRCLK_dly,
	RefSignalName => "CPMDCRCLK",
	RefDelay => ticd_CPMDCRCLK,
	SetupHigh => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(31),
	SetupLow => tsetup_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(31),
	HoldLow => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_posedge_posedge(31),
	HoldHigh => thold_DCRPPCDSDBUSOUT_CPMDCRCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_DCRPPCDSREAD_CPMDCRCLK_posedge,
	TimingData     => Tmkr_DCRPPCDSREAD_CPMDCRCLK_posedge,
	TestSignal     => DCRPPCDSREAD,
	TestSignalName => "DCRPPCDSREAD",
	TestDelay      => 0 ps,
	RefSignal => CPMDCRCLK_dly,
	RefSignalName  => "CPMDCRCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_DCRPPCDSREAD_CPMDCRCLK_posedge_posedge,
	SetupLow       => tsetup_DCRPPCDSREAD_CPMDCRCLK_negedge_posedge,
	HoldLow        => thold_DCRPPCDSREAD_CPMDCRCLK_posedge_posedge,
	HoldHigh       => thold_DCRPPCDSREAD_CPMDCRCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_DCRPPCDSWRITE_CPMDCRCLK_posedge,
	TimingData     => Tmkr_DCRPPCDSWRITE_CPMDCRCLK_posedge,
	TestSignal     => DCRPPCDSWRITE,
	TestSignalName => "DCRPPCDSWRITE",
	TestDelay      => 0 ps,
	RefSignal => CPMDCRCLK_dly,
	RefSignalName  => "CPMDCRCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_DCRPPCDSWRITE_CPMDCRCLK_posedge_posedge,
	SetupLow       => tsetup_DCRPPCDSWRITE_CPMDCRCLK_negedge_posedge,
	HoldLow        => thold_DCRPPCDSWRITE_CPMDCRCLK_posedge_posedge,
	HoldHigh       => thold_DCRPPCDSWRITE_CPMDCRCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_FCMAPUCONFIRMINSTR_CPMFCMCLK_posedge,
	TimingData     => Tmkr_FCMAPUCONFIRMINSTR_CPMFCMCLK_posedge,
	TestSignal     => FCMAPUCONFIRMINSTR,
	TestSignalName => "FCMAPUCONFIRMINSTR",
	TestDelay      => 0 ps,
	RefSignal => CPMFCMCLK_dly,
	RefSignalName  => "CPMFCMCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_FCMAPUCONFIRMINSTR_CPMFCMCLK_posedge_posedge,
	SetupLow       => tsetup_FCMAPUCONFIRMINSTR_CPMFCMCLK_negedge_posedge,
	HoldLow        => thold_FCMAPUCONFIRMINSTR_CPMFCMCLK_posedge_posedge,
	HoldHigh       => thold_FCMAPUCONFIRMINSTR_CPMFCMCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUCR0_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUCR0_CPMFCMCLK_posedge,
	TestSignal => FCMAPUCR_dly(0),
	TestSignalName => "FCMAPUCR(0)",
	TestDelay => tisd_FCMAPUCR_CPMFCMCLK(0),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUCR_CPMFCMCLK_posedge_posedge(0),
	SetupLow => tsetup_FCMAPUCR_CPMFCMCLK_negedge_posedge(0),
	HoldLow => thold_FCMAPUCR_CPMFCMCLK_posedge_posedge(0),
	HoldHigh => thold_FCMAPUCR_CPMFCMCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUCR1_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUCR1_CPMFCMCLK_posedge,
	TestSignal => FCMAPUCR_dly(1),
	TestSignalName => "FCMAPUCR(1)",
	TestDelay => tisd_FCMAPUCR_CPMFCMCLK(1),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUCR_CPMFCMCLK_posedge_posedge(1),
	SetupLow => tsetup_FCMAPUCR_CPMFCMCLK_negedge_posedge(1),
	HoldLow => thold_FCMAPUCR_CPMFCMCLK_posedge_posedge(1),
	HoldHigh => thold_FCMAPUCR_CPMFCMCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUCR2_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUCR2_CPMFCMCLK_posedge,
	TestSignal => FCMAPUCR_dly(2),
	TestSignalName => "FCMAPUCR(2)",
	TestDelay => tisd_FCMAPUCR_CPMFCMCLK(2),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUCR_CPMFCMCLK_posedge_posedge(2),
	SetupLow => tsetup_FCMAPUCR_CPMFCMCLK_negedge_posedge(2),
	HoldLow => thold_FCMAPUCR_CPMFCMCLK_posedge_posedge(2),
	HoldHigh => thold_FCMAPUCR_CPMFCMCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUCR3_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUCR3_CPMFCMCLK_posedge,
	TestSignal => FCMAPUCR_dly(3),
	TestSignalName => "FCMAPUCR(3)",
	TestDelay => tisd_FCMAPUCR_CPMFCMCLK(3),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUCR_CPMFCMCLK_posedge_posedge(3),
	SetupLow => tsetup_FCMAPUCR_CPMFCMCLK_negedge_posedge(3),
	HoldLow => thold_FCMAPUCR_CPMFCMCLK_posedge_posedge(3),
	HoldHigh => thold_FCMAPUCR_CPMFCMCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_FCMAPUDONE_CPMFCMCLK_posedge,
	TimingData     => Tmkr_FCMAPUDONE_CPMFCMCLK_posedge,
	TestSignal     => FCMAPUDONE,
	TestSignalName => "FCMAPUDONE",
	TestDelay      => 0 ps,
	RefSignal => CPMFCMCLK_dly,
	RefSignalName  => "CPMFCMCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_FCMAPUDONE_CPMFCMCLK_posedge_posedge,
	SetupLow       => tsetup_FCMAPUDONE_CPMFCMCLK_negedge_posedge,
	HoldLow        => thold_FCMAPUDONE_CPMFCMCLK_posedge_posedge,
	HoldHigh       => thold_FCMAPUDONE_CPMFCMCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_FCMAPUEXCEPTION_CPMFCMCLK_posedge,
	TimingData     => Tmkr_FCMAPUEXCEPTION_CPMFCMCLK_posedge,
	TestSignal     => FCMAPUEXCEPTION,
	TestSignalName => "FCMAPUEXCEPTION",
	TestDelay      => 0 ps,
	RefSignal => CPMFCMCLK_dly,
	RefSignalName  => "CPMFCMCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_FCMAPUEXCEPTION_CPMFCMCLK_posedge_posedge,
	SetupLow       => tsetup_FCMAPUEXCEPTION_CPMFCMCLK_negedge_posedge,
	HoldLow        => thold_FCMAPUEXCEPTION_CPMFCMCLK_posedge_posedge,
	HoldHigh       => thold_FCMAPUEXCEPTION_CPMFCMCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_FCMAPUFPSCRFEX_CPMFCMCLK_posedge,
	TimingData     => Tmkr_FCMAPUFPSCRFEX_CPMFCMCLK_posedge,
	TestSignal     => FCMAPUFPSCRFEX,
	TestSignalName => "FCMAPUFPSCRFEX",
	TestDelay      => 0 ps,
	RefSignal => CPMFCMCLK_dly,
	RefSignalName  => "CPMFCMCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_FCMAPUFPSCRFEX_CPMFCMCLK_posedge_posedge,
	SetupLow       => tsetup_FCMAPUFPSCRFEX_CPMFCMCLK_negedge_posedge,
	HoldLow        => thold_FCMAPUFPSCRFEX_CPMFCMCLK_posedge_posedge,
	HoldHigh       => thold_FCMAPUFPSCRFEX_CPMFCMCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT0_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT0_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(0),
	TestSignalName => "FCMAPURESULT(0)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(0),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(0),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(0),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(0),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT1_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT1_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(1),
	TestSignalName => "FCMAPURESULT(1)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(1),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(1),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(1),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(1),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT2_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT2_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(2),
	TestSignalName => "FCMAPURESULT(2)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(2),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(2),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(2),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(2),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT3_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT3_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(3),
	TestSignalName => "FCMAPURESULT(3)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(3),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(3),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(3),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(3),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT4_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT4_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(4),
	TestSignalName => "FCMAPURESULT(4)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(4),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(4),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(4),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(4),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT5_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT5_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(5),
	TestSignalName => "FCMAPURESULT(5)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(5),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(5),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(5),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(5),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT6_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT6_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(6),
	TestSignalName => "FCMAPURESULT(6)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(6),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(6),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(6),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(6),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT7_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT7_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(7),
	TestSignalName => "FCMAPURESULT(7)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(7),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(7),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(7),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(7),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT8_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT8_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(8),
	TestSignalName => "FCMAPURESULT(8)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(8),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(8),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(8),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(8),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT9_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT9_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(9),
	TestSignalName => "FCMAPURESULT(9)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(9),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(9),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(9),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(9),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT10_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT10_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(10),
	TestSignalName => "FCMAPURESULT(10)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(10),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(10),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(10),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(10),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT11_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT11_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(11),
	TestSignalName => "FCMAPURESULT(11)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(11),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(11),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(11),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(11),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT12_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT12_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(12),
	TestSignalName => "FCMAPURESULT(12)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(12),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(12),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(12),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(12),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT13_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT13_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(13),
	TestSignalName => "FCMAPURESULT(13)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(13),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(13),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(13),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(13),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT14_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT14_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(14),
	TestSignalName => "FCMAPURESULT(14)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(14),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(14),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(14),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(14),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT15_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT15_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(15),
	TestSignalName => "FCMAPURESULT(15)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(15),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(15),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(15),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(15),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT16_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT16_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(16),
	TestSignalName => "FCMAPURESULT(16)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(16),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(16),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(16),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(16),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(16),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT17_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT17_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(17),
	TestSignalName => "FCMAPURESULT(17)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(17),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(17),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(17),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(17),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(17),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT18_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT18_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(18),
	TestSignalName => "FCMAPURESULT(18)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(18),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(18),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(18),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(18),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(18),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT19_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT19_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(19),
	TestSignalName => "FCMAPURESULT(19)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(19),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(19),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(19),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(19),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(19),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT20_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT20_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(20),
	TestSignalName => "FCMAPURESULT(20)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(20),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(20),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(20),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(20),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(20),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT21_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT21_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(21),
	TestSignalName => "FCMAPURESULT(21)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(21),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(21),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(21),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(21),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(21),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT22_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT22_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(22),
	TestSignalName => "FCMAPURESULT(22)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(22),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(22),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(22),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(22),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(22),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT23_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT23_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(23),
	TestSignalName => "FCMAPURESULT(23)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(23),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(23),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(23),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(23),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(23),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT24_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT24_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(24),
	TestSignalName => "FCMAPURESULT(24)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(24),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(24),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(24),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(24),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(24),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT25_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT25_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(25),
	TestSignalName => "FCMAPURESULT(25)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(25),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(25),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(25),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(25),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(25),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT26_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT26_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(26),
	TestSignalName => "FCMAPURESULT(26)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(26),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(26),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(26),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(26),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(26),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT27_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT27_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(27),
	TestSignalName => "FCMAPURESULT(27)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(27),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(27),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(27),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(27),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(27),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT28_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT28_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(28),
	TestSignalName => "FCMAPURESULT(28)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(28),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(28),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(28),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(28),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT29_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT29_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(29),
	TestSignalName => "FCMAPURESULT(29)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(29),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(29),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(29),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(29),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT30_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT30_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(30),
	TestSignalName => "FCMAPURESULT(30)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(30),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(30),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(30),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(30),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPURESULT31_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPURESULT31_CPMFCMCLK_posedge,
	TestSignal => FCMAPURESULT_dly(31),
	TestSignalName => "FCMAPURESULT(31)",
	TestDelay => tisd_FCMAPURESULT_CPMFCMCLK(31),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPURESULT_CPMFCMCLK_posedge_posedge(31),
	SetupLow => tsetup_FCMAPURESULT_CPMFCMCLK_negedge_posedge(31),
	HoldLow => thold_FCMAPURESULT_CPMFCMCLK_posedge_posedge(31),
	HoldHigh => thold_FCMAPURESULT_CPMFCMCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_FCMAPURESULTVALID_CPMFCMCLK_posedge,
	TimingData     => Tmkr_FCMAPURESULTVALID_CPMFCMCLK_posedge,
	TestSignal     => FCMAPURESULTVALID,
	TestSignalName => "FCMAPURESULTVALID",
	TestDelay      => 0 ps,
	RefSignal => CPMFCMCLK_dly,
	RefSignalName  => "CPMFCMCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_FCMAPURESULTVALID_CPMFCMCLK_posedge_posedge,
	SetupLow       => tsetup_FCMAPURESULTVALID_CPMFCMCLK_negedge_posedge,
	HoldLow        => thold_FCMAPURESULTVALID_CPMFCMCLK_posedge_posedge,
	HoldHigh       => thold_FCMAPURESULTVALID_CPMFCMCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_FCMAPUSLEEPNOTREADY_CPMFCMCLK_posedge,
	TimingData     => Tmkr_FCMAPUSLEEPNOTREADY_CPMFCMCLK_posedge,
	TestSignal     => FCMAPUSLEEPNOTREADY,
	TestSignalName => "FCMAPUSLEEPNOTREADY",
	TestDelay      => 0 ps,
	RefSignal => CPMFCMCLK_dly,
	RefSignalName  => "CPMFCMCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_FCMAPUSLEEPNOTREADY_CPMFCMCLK_posedge_posedge,
	SetupLow       => tsetup_FCMAPUSLEEPNOTREADY_CPMFCMCLK_negedge_posedge,
	HoldLow        => thold_FCMAPUSLEEPNOTREADY_CPMFCMCLK_posedge_posedge,
	HoldHigh       => thold_FCMAPUSLEEPNOTREADY_CPMFCMCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA0_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA0_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(0),
	TestSignalName => "FCMAPUSTOREDATA(0)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(0),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(0),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(0),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(0),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA1_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA1_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(1),
	TestSignalName => "FCMAPUSTOREDATA(1)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(1),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(1),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(1),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(1),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA2_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA2_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(2),
	TestSignalName => "FCMAPUSTOREDATA(2)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(2),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(2),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(2),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(2),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA3_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA3_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(3),
	TestSignalName => "FCMAPUSTOREDATA(3)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(3),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(3),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(3),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(3),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA4_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA4_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(4),
	TestSignalName => "FCMAPUSTOREDATA(4)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(4),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(4),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(4),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(4),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA5_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA5_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(5),
	TestSignalName => "FCMAPUSTOREDATA(5)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(5),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(5),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(5),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(5),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA6_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA6_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(6),
	TestSignalName => "FCMAPUSTOREDATA(6)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(6),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(6),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(6),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(6),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA7_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA7_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(7),
	TestSignalName => "FCMAPUSTOREDATA(7)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(7),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(7),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(7),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(7),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA8_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA8_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(8),
	TestSignalName => "FCMAPUSTOREDATA(8)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(8),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(8),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(8),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(8),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA9_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA9_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(9),
	TestSignalName => "FCMAPUSTOREDATA(9)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(9),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(9),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(9),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(9),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA10_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA10_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(10),
	TestSignalName => "FCMAPUSTOREDATA(10)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(10),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(10),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(10),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(10),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA11_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA11_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(11),
	TestSignalName => "FCMAPUSTOREDATA(11)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(11),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(11),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(11),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(11),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA12_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA12_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(12),
	TestSignalName => "FCMAPUSTOREDATA(12)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(12),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(12),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(12),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(12),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA13_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA13_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(13),
	TestSignalName => "FCMAPUSTOREDATA(13)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(13),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(13),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(13),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(13),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA14_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA14_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(14),
	TestSignalName => "FCMAPUSTOREDATA(14)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(14),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(14),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(14),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(14),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA15_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA15_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(15),
	TestSignalName => "FCMAPUSTOREDATA(15)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(15),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(15),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(15),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(15),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA16_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA16_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(16),
	TestSignalName => "FCMAPUSTOREDATA(16)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(16),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(16),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(16),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(16),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(16),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA17_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA17_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(17),
	TestSignalName => "FCMAPUSTOREDATA(17)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(17),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(17),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(17),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(17),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(17),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA18_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA18_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(18),
	TestSignalName => "FCMAPUSTOREDATA(18)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(18),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(18),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(18),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(18),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(18),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA19_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA19_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(19),
	TestSignalName => "FCMAPUSTOREDATA(19)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(19),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(19),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(19),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(19),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(19),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA20_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA20_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(20),
	TestSignalName => "FCMAPUSTOREDATA(20)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(20),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(20),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(20),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(20),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(20),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA21_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA21_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(21),
	TestSignalName => "FCMAPUSTOREDATA(21)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(21),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(21),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(21),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(21),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(21),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA22_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA22_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(22),
	TestSignalName => "FCMAPUSTOREDATA(22)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(22),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(22),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(22),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(22),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(22),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA23_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA23_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(23),
	TestSignalName => "FCMAPUSTOREDATA(23)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(23),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(23),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(23),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(23),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(23),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA24_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA24_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(24),
	TestSignalName => "FCMAPUSTOREDATA(24)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(24),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(24),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(24),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(24),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(24),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA25_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA25_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(25),
	TestSignalName => "FCMAPUSTOREDATA(25)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(25),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(25),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(25),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(25),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(25),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA26_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA26_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(26),
	TestSignalName => "FCMAPUSTOREDATA(26)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(26),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(26),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(26),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(26),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(26),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA27_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA27_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(27),
	TestSignalName => "FCMAPUSTOREDATA(27)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(27),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(27),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(27),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(27),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(27),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA28_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA28_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(28),
	TestSignalName => "FCMAPUSTOREDATA(28)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(28),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(28),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(28),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(28),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA29_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA29_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(29),
	TestSignalName => "FCMAPUSTOREDATA(29)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(29),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(29),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(29),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(29),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA30_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA30_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(30),
	TestSignalName => "FCMAPUSTOREDATA(30)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(30),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(30),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(30),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(30),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA31_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA31_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(31),
	TestSignalName => "FCMAPUSTOREDATA(31)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(31),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(31),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(31),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(31),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA32_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA32_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(32),
	TestSignalName => "FCMAPUSTOREDATA(32)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(32),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(32),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(32),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(32),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(32),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA33_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA33_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(33),
	TestSignalName => "FCMAPUSTOREDATA(33)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(33),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(33),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(33),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(33),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(33),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA34_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA34_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(34),
	TestSignalName => "FCMAPUSTOREDATA(34)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(34),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(34),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(34),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(34),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(34),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA35_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA35_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(35),
	TestSignalName => "FCMAPUSTOREDATA(35)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(35),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(35),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(35),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(35),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(35),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA36_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA36_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(36),
	TestSignalName => "FCMAPUSTOREDATA(36)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(36),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(36),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(36),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(36),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(36),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA37_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA37_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(37),
	TestSignalName => "FCMAPUSTOREDATA(37)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(37),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(37),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(37),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(37),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(37),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA38_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA38_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(38),
	TestSignalName => "FCMAPUSTOREDATA(38)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(38),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(38),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(38),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(38),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(38),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA39_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA39_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(39),
	TestSignalName => "FCMAPUSTOREDATA(39)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(39),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(39),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(39),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(39),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(39),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA40_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA40_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(40),
	TestSignalName => "FCMAPUSTOREDATA(40)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(40),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(40),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(40),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(40),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(40),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA41_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA41_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(41),
	TestSignalName => "FCMAPUSTOREDATA(41)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(41),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(41),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(41),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(41),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(41),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA42_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA42_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(42),
	TestSignalName => "FCMAPUSTOREDATA(42)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(42),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(42),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(42),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(42),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(42),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA43_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA43_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(43),
	TestSignalName => "FCMAPUSTOREDATA(43)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(43),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(43),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(43),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(43),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(43),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA44_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA44_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(44),
	TestSignalName => "FCMAPUSTOREDATA(44)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(44),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(44),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(44),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(44),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(44),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA45_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA45_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(45),
	TestSignalName => "FCMAPUSTOREDATA(45)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(45),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(45),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(45),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(45),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(45),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA46_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA46_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(46),
	TestSignalName => "FCMAPUSTOREDATA(46)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(46),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(46),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(46),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(46),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(46),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA47_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA47_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(47),
	TestSignalName => "FCMAPUSTOREDATA(47)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(47),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(47),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(47),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(47),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(47),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA48_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA48_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(48),
	TestSignalName => "FCMAPUSTOREDATA(48)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(48),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(48),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(48),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(48),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(48),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA49_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA49_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(49),
	TestSignalName => "FCMAPUSTOREDATA(49)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(49),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(49),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(49),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(49),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(49),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA50_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA50_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(50),
	TestSignalName => "FCMAPUSTOREDATA(50)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(50),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(50),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(50),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(50),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(50),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA51_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA51_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(51),
	TestSignalName => "FCMAPUSTOREDATA(51)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(51),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(51),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(51),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(51),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(51),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA52_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA52_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(52),
	TestSignalName => "FCMAPUSTOREDATA(52)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(52),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(52),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(52),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(52),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(52),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA53_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA53_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(53),
	TestSignalName => "FCMAPUSTOREDATA(53)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(53),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(53),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(53),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(53),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(53),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA54_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA54_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(54),
	TestSignalName => "FCMAPUSTOREDATA(54)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(54),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(54),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(54),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(54),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(54),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA55_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA55_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(55),
	TestSignalName => "FCMAPUSTOREDATA(55)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(55),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(55),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(55),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(55),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(55),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA56_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA56_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(56),
	TestSignalName => "FCMAPUSTOREDATA(56)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(56),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(56),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(56),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(56),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(56),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA57_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA57_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(57),
	TestSignalName => "FCMAPUSTOREDATA(57)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(57),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(57),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(57),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(57),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(57),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA58_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA58_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(58),
	TestSignalName => "FCMAPUSTOREDATA(58)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(58),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(58),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(58),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(58),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(58),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA59_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA59_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(59),
	TestSignalName => "FCMAPUSTOREDATA(59)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(59),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(59),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(59),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(59),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(59),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA60_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA60_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(60),
	TestSignalName => "FCMAPUSTOREDATA(60)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(60),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(60),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(60),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(60),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(60),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA61_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA61_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(61),
	TestSignalName => "FCMAPUSTOREDATA(61)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(61),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(61),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(61),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(61),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(61),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA62_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA62_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(62),
	TestSignalName => "FCMAPUSTOREDATA(62)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(62),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(62),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(62),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(62),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(62),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA63_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA63_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(63),
	TestSignalName => "FCMAPUSTOREDATA(63)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(63),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(63),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(63),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(63),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(63),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA64_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA64_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(64),
	TestSignalName => "FCMAPUSTOREDATA(64)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(64),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(64),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(64),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(64),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(64),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA65_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA65_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(65),
	TestSignalName => "FCMAPUSTOREDATA(65)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(65),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(65),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(65),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(65),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(65),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA66_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA66_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(66),
	TestSignalName => "FCMAPUSTOREDATA(66)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(66),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(66),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(66),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(66),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(66),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA67_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA67_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(67),
	TestSignalName => "FCMAPUSTOREDATA(67)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(67),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(67),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(67),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(67),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(67),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA68_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA68_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(68),
	TestSignalName => "FCMAPUSTOREDATA(68)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(68),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(68),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(68),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(68),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(68),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA69_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA69_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(69),
	TestSignalName => "FCMAPUSTOREDATA(69)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(69),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(69),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(69),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(69),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(69),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA70_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA70_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(70),
	TestSignalName => "FCMAPUSTOREDATA(70)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(70),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(70),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(70),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(70),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(70),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA71_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA71_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(71),
	TestSignalName => "FCMAPUSTOREDATA(71)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(71),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(71),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(71),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(71),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(71),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA72_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA72_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(72),
	TestSignalName => "FCMAPUSTOREDATA(72)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(72),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(72),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(72),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(72),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(72),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA73_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA73_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(73),
	TestSignalName => "FCMAPUSTOREDATA(73)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(73),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(73),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(73),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(73),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(73),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA74_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA74_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(74),
	TestSignalName => "FCMAPUSTOREDATA(74)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(74),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(74),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(74),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(74),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(74),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA75_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA75_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(75),
	TestSignalName => "FCMAPUSTOREDATA(75)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(75),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(75),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(75),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(75),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(75),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA76_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA76_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(76),
	TestSignalName => "FCMAPUSTOREDATA(76)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(76),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(76),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(76),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(76),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(76),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA77_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA77_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(77),
	TestSignalName => "FCMAPUSTOREDATA(77)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(77),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(77),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(77),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(77),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(77),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA78_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA78_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(78),
	TestSignalName => "FCMAPUSTOREDATA(78)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(78),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(78),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(78),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(78),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(78),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA79_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA79_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(79),
	TestSignalName => "FCMAPUSTOREDATA(79)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(79),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(79),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(79),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(79),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(79),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA80_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA80_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(80),
	TestSignalName => "FCMAPUSTOREDATA(80)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(80),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(80),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(80),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(80),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(80),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA81_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA81_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(81),
	TestSignalName => "FCMAPUSTOREDATA(81)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(81),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(81),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(81),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(81),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(81),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA82_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA82_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(82),
	TestSignalName => "FCMAPUSTOREDATA(82)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(82),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(82),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(82),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(82),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(82),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA83_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA83_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(83),
	TestSignalName => "FCMAPUSTOREDATA(83)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(83),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(83),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(83),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(83),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(83),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA84_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA84_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(84),
	TestSignalName => "FCMAPUSTOREDATA(84)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(84),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(84),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(84),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(84),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(84),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA85_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA85_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(85),
	TestSignalName => "FCMAPUSTOREDATA(85)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(85),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(85),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(85),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(85),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(85),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA86_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA86_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(86),
	TestSignalName => "FCMAPUSTOREDATA(86)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(86),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(86),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(86),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(86),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(86),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA87_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA87_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(87),
	TestSignalName => "FCMAPUSTOREDATA(87)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(87),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(87),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(87),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(87),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(87),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA88_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA88_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(88),
	TestSignalName => "FCMAPUSTOREDATA(88)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(88),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(88),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(88),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(88),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(88),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA89_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA89_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(89),
	TestSignalName => "FCMAPUSTOREDATA(89)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(89),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(89),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(89),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(89),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(89),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA90_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA90_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(90),
	TestSignalName => "FCMAPUSTOREDATA(90)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(90),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(90),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(90),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(90),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(90),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA91_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA91_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(91),
	TestSignalName => "FCMAPUSTOREDATA(91)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(91),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(91),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(91),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(91),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(91),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA92_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA92_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(92),
	TestSignalName => "FCMAPUSTOREDATA(92)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(92),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(92),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(92),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(92),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(92),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA93_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA93_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(93),
	TestSignalName => "FCMAPUSTOREDATA(93)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(93),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(93),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(93),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(93),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(93),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA94_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA94_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(94),
	TestSignalName => "FCMAPUSTOREDATA(94)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(94),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(94),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(94),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(94),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(94),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA95_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA95_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(95),
	TestSignalName => "FCMAPUSTOREDATA(95)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(95),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(95),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(95),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(95),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(95),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA96_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA96_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(96),
	TestSignalName => "FCMAPUSTOREDATA(96)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(96),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(96),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(96),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(96),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(96),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA97_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA97_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(97),
	TestSignalName => "FCMAPUSTOREDATA(97)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(97),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(97),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(97),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(97),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(97),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA98_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA98_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(98),
	TestSignalName => "FCMAPUSTOREDATA(98)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(98),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(98),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(98),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(98),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(98),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA99_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA99_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(99),
	TestSignalName => "FCMAPUSTOREDATA(99)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(99),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(99),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(99),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(99),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(99),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA100_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA100_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(100),
	TestSignalName => "FCMAPUSTOREDATA(100)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(100),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(100),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(100),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(100),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(100),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA101_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA101_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(101),
	TestSignalName => "FCMAPUSTOREDATA(101)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(101),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(101),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(101),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(101),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(101),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA102_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA102_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(102),
	TestSignalName => "FCMAPUSTOREDATA(102)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(102),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(102),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(102),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(102),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(102),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA103_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA103_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(103),
	TestSignalName => "FCMAPUSTOREDATA(103)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(103),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(103),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(103),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(103),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(103),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA104_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA104_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(104),
	TestSignalName => "FCMAPUSTOREDATA(104)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(104),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(104),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(104),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(104),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(104),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA105_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA105_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(105),
	TestSignalName => "FCMAPUSTOREDATA(105)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(105),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(105),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(105),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(105),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(105),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA106_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA106_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(106),
	TestSignalName => "FCMAPUSTOREDATA(106)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(106),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(106),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(106),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(106),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(106),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA107_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA107_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(107),
	TestSignalName => "FCMAPUSTOREDATA(107)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(107),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(107),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(107),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(107),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(107),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA108_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA108_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(108),
	TestSignalName => "FCMAPUSTOREDATA(108)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(108),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(108),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(108),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(108),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(108),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA109_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA109_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(109),
	TestSignalName => "FCMAPUSTOREDATA(109)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(109),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(109),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(109),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(109),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(109),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA110_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA110_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(110),
	TestSignalName => "FCMAPUSTOREDATA(110)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(110),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(110),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(110),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(110),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(110),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA111_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA111_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(111),
	TestSignalName => "FCMAPUSTOREDATA(111)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(111),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(111),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(111),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(111),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(111),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA112_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA112_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(112),
	TestSignalName => "FCMAPUSTOREDATA(112)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(112),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(112),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(112),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(112),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(112),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA113_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA113_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(113),
	TestSignalName => "FCMAPUSTOREDATA(113)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(113),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(113),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(113),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(113),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(113),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA114_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA114_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(114),
	TestSignalName => "FCMAPUSTOREDATA(114)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(114),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(114),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(114),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(114),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(114),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA115_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA115_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(115),
	TestSignalName => "FCMAPUSTOREDATA(115)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(115),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(115),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(115),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(115),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(115),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA116_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA116_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(116),
	TestSignalName => "FCMAPUSTOREDATA(116)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(116),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(116),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(116),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(116),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(116),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA117_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA117_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(117),
	TestSignalName => "FCMAPUSTOREDATA(117)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(117),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(117),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(117),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(117),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(117),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA118_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA118_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(118),
	TestSignalName => "FCMAPUSTOREDATA(118)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(118),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(118),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(118),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(118),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(118),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA119_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA119_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(119),
	TestSignalName => "FCMAPUSTOREDATA(119)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(119),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(119),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(119),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(119),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(119),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA120_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA120_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(120),
	TestSignalName => "FCMAPUSTOREDATA(120)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(120),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(120),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(120),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(120),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(120),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA121_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA121_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(121),
	TestSignalName => "FCMAPUSTOREDATA(121)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(121),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(121),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(121),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(121),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(121),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA122_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA122_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(122),
	TestSignalName => "FCMAPUSTOREDATA(122)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(122),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(122),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(122),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(122),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(122),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA123_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA123_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(123),
	TestSignalName => "FCMAPUSTOREDATA(123)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(123),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(123),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(123),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(123),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(123),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA124_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA124_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(124),
	TestSignalName => "FCMAPUSTOREDATA(124)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(124),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(124),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(124),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(124),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(124),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA125_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA125_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(125),
	TestSignalName => "FCMAPUSTOREDATA(125)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(125),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(125),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(125),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(125),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(125),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA126_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA126_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(126),
	TestSignalName => "FCMAPUSTOREDATA(126)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(126),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(126),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(126),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(126),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(126),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_FCMAPUSTOREDATA127_CPMFCMCLK_posedge,
	TimingData => Tmkr_FCMAPUSTOREDATA127_CPMFCMCLK_posedge,
	TestSignal => FCMAPUSTOREDATA_dly(127),
	TestSignalName => "FCMAPUSTOREDATA(127)",
	TestDelay => tisd_FCMAPUSTOREDATA_CPMFCMCLK(127),
	RefSignal => CPMFCMCLK_dly,
	RefSignalName => "CPMFCMCLK",
	RefDelay => ticd_CPMFCMCLK,
	SetupHigh => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(127),
	SetupLow => tsetup_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(127),
	HoldLow => thold_FCMAPUSTOREDATA_CPMFCMCLK_posedge_posedge(127),
	HoldHigh => thold_FCMAPUSTOREDATA_CPMFCMCLK_negedge_posedge(127),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_JTGC440TDI_JTGC440TCK_posedge,
	TimingData     => Tmkr_JTGC440TDI_JTGC440TCK_posedge,
	TestSignal     => JTGC440TDI,
	TestSignalName => "JTGC440TDI",
	TestDelay      => 0 ps,
	RefSignal => JTGC440TCK_dly,
	RefSignalName  => "JTGC440TCK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_JTGC440TDI_JTGC440TCK_posedge_posedge,
	SetupLow       => tsetup_JTGC440TDI_JTGC440TCK_negedge_posedge,
	HoldLow        => thold_JTGC440TDI_JTGC440TCK_posedge_posedge,
	HoldHigh       => thold_JTGC440TDI_JTGC440TCK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_JTGC440TMS_JTGC440TCK_posedge,
	TimingData     => Tmkr_JTGC440TMS_JTGC440TCK_posedge,
	TestSignal     => JTGC440TMS,
	TestSignalName => "JTGC440TMS",
	TestDelay      => 0 ps,
	RefSignal => JTGC440TCK_dly,
	RefSignalName  => "JTGC440TCK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_JTGC440TMS_JTGC440TCK_posedge_posedge,
	SetupLow       => tsetup_JTGC440TMS_JTGC440TCK_negedge_posedge,
	HoldLow        => thold_JTGC440TMS_JTGC440TCK_posedge_posedge,
	HoldHigh       => thold_JTGC440TMS_JTGC440TCK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_MCMIADDRREADYTOACCEPT_CPMMCCLK_posedge,
	TimingData     => Tmkr_MCMIADDRREADYTOACCEPT_CPMMCCLK_posedge,
	TestSignal     => MCMIADDRREADYTOACCEPT,
	TestSignalName => "MCMIADDRREADYTOACCEPT",
	TestDelay      => 0 ps,
	RefSignal => CPMMCCLK_dly,
	RefSignalName  => "CPMMCCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_MCMIADDRREADYTOACCEPT_CPMMCCLK_posedge_posedge,
	SetupLow       => tsetup_MCMIADDRREADYTOACCEPT_CPMMCCLK_negedge_posedge,
	HoldLow        => thold_MCMIADDRREADYTOACCEPT_CPMMCCLK_posedge_posedge,
	HoldHigh       => thold_MCMIADDRREADYTOACCEPT_CPMMCCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA0_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA0_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(0),
	TestSignalName => "MCMIREADDATA(0)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(0),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(0),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(0),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(0),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(0),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA1_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA1_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(1),
	TestSignalName => "MCMIREADDATA(1)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(1),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(1),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(1),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(1),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(1),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA2_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA2_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(2),
	TestSignalName => "MCMIREADDATA(2)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(2),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(2),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(2),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(2),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(2),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA3_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA3_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(3),
	TestSignalName => "MCMIREADDATA(3)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(3),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(3),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(3),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(3),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(3),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA4_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA4_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(4),
	TestSignalName => "MCMIREADDATA(4)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(4),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(4),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(4),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(4),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(4),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA5_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA5_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(5),
	TestSignalName => "MCMIREADDATA(5)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(5),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(5),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(5),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(5),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(5),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA6_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA6_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(6),
	TestSignalName => "MCMIREADDATA(6)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(6),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(6),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(6),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(6),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(6),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA7_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA7_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(7),
	TestSignalName => "MCMIREADDATA(7)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(7),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(7),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(7),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(7),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(7),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA8_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA8_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(8),
	TestSignalName => "MCMIREADDATA(8)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(8),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(8),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(8),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(8),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(8),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA9_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA9_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(9),
	TestSignalName => "MCMIREADDATA(9)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(9),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(9),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(9),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(9),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(9),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA10_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA10_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(10),
	TestSignalName => "MCMIREADDATA(10)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(10),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(10),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(10),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(10),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(10),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA11_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA11_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(11),
	TestSignalName => "MCMIREADDATA(11)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(11),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(11),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(11),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(11),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(11),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA12_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA12_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(12),
	TestSignalName => "MCMIREADDATA(12)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(12),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(12),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(12),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(12),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(12),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA13_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA13_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(13),
	TestSignalName => "MCMIREADDATA(13)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(13),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(13),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(13),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(13),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(13),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA14_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA14_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(14),
	TestSignalName => "MCMIREADDATA(14)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(14),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(14),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(14),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(14),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(14),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA15_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA15_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(15),
	TestSignalName => "MCMIREADDATA(15)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(15),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(15),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(15),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(15),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(15),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA16_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA16_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(16),
	TestSignalName => "MCMIREADDATA(16)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(16),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(16),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(16),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(16),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(16),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA17_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA17_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(17),
	TestSignalName => "MCMIREADDATA(17)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(17),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(17),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(17),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(17),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(17),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA18_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA18_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(18),
	TestSignalName => "MCMIREADDATA(18)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(18),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(18),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(18),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(18),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(18),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA19_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA19_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(19),
	TestSignalName => "MCMIREADDATA(19)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(19),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(19),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(19),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(19),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(19),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA20_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA20_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(20),
	TestSignalName => "MCMIREADDATA(20)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(20),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(20),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(20),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(20),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(20),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA21_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA21_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(21),
	TestSignalName => "MCMIREADDATA(21)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(21),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(21),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(21),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(21),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(21),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA22_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA22_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(22),
	TestSignalName => "MCMIREADDATA(22)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(22),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(22),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(22),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(22),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(22),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA23_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA23_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(23),
	TestSignalName => "MCMIREADDATA(23)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(23),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(23),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(23),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(23),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(23),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA24_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA24_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(24),
	TestSignalName => "MCMIREADDATA(24)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(24),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(24),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(24),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(24),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(24),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA25_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA25_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(25),
	TestSignalName => "MCMIREADDATA(25)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(25),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(25),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(25),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(25),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(25),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA26_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA26_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(26),
	TestSignalName => "MCMIREADDATA(26)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(26),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(26),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(26),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(26),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(26),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA27_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA27_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(27),
	TestSignalName => "MCMIREADDATA(27)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(27),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(27),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(27),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(27),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(27),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA28_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA28_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(28),
	TestSignalName => "MCMIREADDATA(28)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(28),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(28),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(28),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(28),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(28),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA29_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA29_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(29),
	TestSignalName => "MCMIREADDATA(29)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(29),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(29),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(29),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(29),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(29),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA30_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA30_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(30),
	TestSignalName => "MCMIREADDATA(30)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(30),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(30),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(30),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(30),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(30),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA31_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA31_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(31),
	TestSignalName => "MCMIREADDATA(31)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(31),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(31),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(31),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(31),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(31),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA32_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA32_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(32),
	TestSignalName => "MCMIREADDATA(32)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(32),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(32),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(32),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(32),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(32),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA33_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA33_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(33),
	TestSignalName => "MCMIREADDATA(33)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(33),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(33),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(33),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(33),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(33),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA34_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA34_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(34),
	TestSignalName => "MCMIREADDATA(34)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(34),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(34),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(34),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(34),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(34),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA35_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA35_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(35),
	TestSignalName => "MCMIREADDATA(35)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(35),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(35),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(35),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(35),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(35),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA36_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA36_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(36),
	TestSignalName => "MCMIREADDATA(36)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(36),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(36),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(36),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(36),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(36),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA37_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA37_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(37),
	TestSignalName => "MCMIREADDATA(37)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(37),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(37),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(37),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(37),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(37),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA38_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA38_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(38),
	TestSignalName => "MCMIREADDATA(38)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(38),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(38),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(38),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(38),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(38),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA39_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA39_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(39),
	TestSignalName => "MCMIREADDATA(39)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(39),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(39),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(39),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(39),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(39),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA40_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA40_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(40),
	TestSignalName => "MCMIREADDATA(40)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(40),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(40),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(40),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(40),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(40),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA41_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA41_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(41),
	TestSignalName => "MCMIREADDATA(41)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(41),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(41),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(41),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(41),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(41),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA42_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA42_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(42),
	TestSignalName => "MCMIREADDATA(42)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(42),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(42),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(42),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(42),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(42),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA43_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA43_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(43),
	TestSignalName => "MCMIREADDATA(43)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(43),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(43),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(43),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(43),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(43),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA44_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA44_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(44),
	TestSignalName => "MCMIREADDATA(44)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(44),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(44),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(44),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(44),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(44),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA45_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA45_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(45),
	TestSignalName => "MCMIREADDATA(45)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(45),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(45),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(45),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(45),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(45),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA46_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA46_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(46),
	TestSignalName => "MCMIREADDATA(46)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(46),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(46),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(46),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(46),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(46),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA47_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA47_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(47),
	TestSignalName => "MCMIREADDATA(47)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(47),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(47),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(47),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(47),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(47),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA48_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA48_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(48),
	TestSignalName => "MCMIREADDATA(48)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(48),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(48),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(48),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(48),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(48),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA49_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA49_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(49),
	TestSignalName => "MCMIREADDATA(49)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(49),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(49),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(49),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(49),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(49),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA50_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA50_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(50),
	TestSignalName => "MCMIREADDATA(50)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(50),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(50),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(50),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(50),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(50),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA51_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA51_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(51),
	TestSignalName => "MCMIREADDATA(51)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(51),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(51),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(51),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(51),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(51),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA52_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA52_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(52),
	TestSignalName => "MCMIREADDATA(52)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(52),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(52),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(52),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(52),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(52),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA53_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA53_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(53),
	TestSignalName => "MCMIREADDATA(53)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(53),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(53),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(53),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(53),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(53),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA54_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA54_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(54),
	TestSignalName => "MCMIREADDATA(54)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(54),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(54),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(54),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(54),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(54),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA55_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA55_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(55),
	TestSignalName => "MCMIREADDATA(55)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(55),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(55),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(55),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(55),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(55),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA56_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA56_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(56),
	TestSignalName => "MCMIREADDATA(56)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(56),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(56),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(56),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(56),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(56),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA57_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA57_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(57),
	TestSignalName => "MCMIREADDATA(57)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(57),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(57),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(57),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(57),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(57),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA58_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA58_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(58),
	TestSignalName => "MCMIREADDATA(58)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(58),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(58),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(58),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(58),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(58),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA59_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA59_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(59),
	TestSignalName => "MCMIREADDATA(59)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(59),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(59),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(59),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(59),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(59),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA60_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA60_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(60),
	TestSignalName => "MCMIREADDATA(60)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(60),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(60),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(60),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(60),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(60),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA61_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA61_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(61),
	TestSignalName => "MCMIREADDATA(61)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(61),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(61),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(61),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(61),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(61),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA62_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA62_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(62),
	TestSignalName => "MCMIREADDATA(62)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(62),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(62),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(62),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(62),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(62),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA63_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA63_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(63),
	TestSignalName => "MCMIREADDATA(63)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(63),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(63),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(63),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(63),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(63),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA64_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA64_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(64),
	TestSignalName => "MCMIREADDATA(64)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(64),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(64),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(64),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(64),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(64),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA65_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA65_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(65),
	TestSignalName => "MCMIREADDATA(65)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(65),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(65),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(65),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(65),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(65),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA66_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA66_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(66),
	TestSignalName => "MCMIREADDATA(66)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(66),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(66),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(66),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(66),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(66),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA67_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA67_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(67),
	TestSignalName => "MCMIREADDATA(67)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(67),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(67),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(67),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(67),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(67),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA68_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA68_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(68),
	TestSignalName => "MCMIREADDATA(68)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(68),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(68),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(68),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(68),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(68),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA69_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA69_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(69),
	TestSignalName => "MCMIREADDATA(69)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(69),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(69),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(69),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(69),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(69),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA70_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA70_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(70),
	TestSignalName => "MCMIREADDATA(70)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(70),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(70),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(70),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(70),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(70),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA71_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA71_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(71),
	TestSignalName => "MCMIREADDATA(71)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(71),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(71),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(71),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(71),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(71),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA72_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA72_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(72),
	TestSignalName => "MCMIREADDATA(72)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(72),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(72),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(72),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(72),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(72),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA73_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA73_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(73),
	TestSignalName => "MCMIREADDATA(73)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(73),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(73),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(73),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(73),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(73),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA74_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA74_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(74),
	TestSignalName => "MCMIREADDATA(74)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(74),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(74),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(74),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(74),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(74),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA75_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA75_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(75),
	TestSignalName => "MCMIREADDATA(75)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(75),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(75),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(75),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(75),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(75),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA76_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA76_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(76),
	TestSignalName => "MCMIREADDATA(76)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(76),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(76),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(76),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(76),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(76),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA77_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA77_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(77),
	TestSignalName => "MCMIREADDATA(77)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(77),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(77),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(77),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(77),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(77),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA78_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA78_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(78),
	TestSignalName => "MCMIREADDATA(78)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(78),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(78),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(78),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(78),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(78),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA79_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA79_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(79),
	TestSignalName => "MCMIREADDATA(79)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(79),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(79),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(79),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(79),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(79),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA80_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA80_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(80),
	TestSignalName => "MCMIREADDATA(80)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(80),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(80),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(80),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(80),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(80),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA81_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA81_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(81),
	TestSignalName => "MCMIREADDATA(81)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(81),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(81),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(81),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(81),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(81),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA82_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA82_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(82),
	TestSignalName => "MCMIREADDATA(82)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(82),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(82),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(82),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(82),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(82),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA83_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA83_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(83),
	TestSignalName => "MCMIREADDATA(83)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(83),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(83),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(83),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(83),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(83),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA84_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA84_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(84),
	TestSignalName => "MCMIREADDATA(84)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(84),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(84),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(84),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(84),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(84),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA85_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA85_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(85),
	TestSignalName => "MCMIREADDATA(85)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(85),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(85),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(85),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(85),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(85),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA86_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA86_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(86),
	TestSignalName => "MCMIREADDATA(86)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(86),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(86),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(86),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(86),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(86),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA87_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA87_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(87),
	TestSignalName => "MCMIREADDATA(87)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(87),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(87),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(87),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(87),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(87),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA88_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA88_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(88),
	TestSignalName => "MCMIREADDATA(88)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(88),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(88),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(88),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(88),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(88),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA89_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA89_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(89),
	TestSignalName => "MCMIREADDATA(89)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(89),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(89),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(89),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(89),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(89),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA90_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA90_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(90),
	TestSignalName => "MCMIREADDATA(90)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(90),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(90),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(90),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(90),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(90),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA91_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA91_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(91),
	TestSignalName => "MCMIREADDATA(91)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(91),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(91),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(91),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(91),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(91),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA92_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA92_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(92),
	TestSignalName => "MCMIREADDATA(92)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(92),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(92),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(92),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(92),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(92),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA93_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA93_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(93),
	TestSignalName => "MCMIREADDATA(93)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(93),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(93),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(93),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(93),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(93),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA94_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA94_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(94),
	TestSignalName => "MCMIREADDATA(94)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(94),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(94),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(94),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(94),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(94),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA95_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA95_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(95),
	TestSignalName => "MCMIREADDATA(95)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(95),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(95),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(95),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(95),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(95),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA96_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA96_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(96),
	TestSignalName => "MCMIREADDATA(96)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(96),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(96),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(96),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(96),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(96),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA97_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA97_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(97),
	TestSignalName => "MCMIREADDATA(97)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(97),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(97),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(97),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(97),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(97),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA98_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA98_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(98),
	TestSignalName => "MCMIREADDATA(98)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(98),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(98),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(98),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(98),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(98),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA99_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA99_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(99),
	TestSignalName => "MCMIREADDATA(99)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(99),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(99),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(99),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(99),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(99),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA100_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA100_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(100),
	TestSignalName => "MCMIREADDATA(100)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(100),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(100),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(100),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(100),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(100),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA101_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA101_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(101),
	TestSignalName => "MCMIREADDATA(101)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(101),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(101),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(101),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(101),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(101),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA102_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA102_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(102),
	TestSignalName => "MCMIREADDATA(102)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(102),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(102),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(102),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(102),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(102),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA103_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA103_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(103),
	TestSignalName => "MCMIREADDATA(103)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(103),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(103),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(103),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(103),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(103),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA104_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA104_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(104),
	TestSignalName => "MCMIREADDATA(104)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(104),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(104),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(104),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(104),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(104),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA105_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA105_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(105),
	TestSignalName => "MCMIREADDATA(105)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(105),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(105),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(105),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(105),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(105),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA106_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA106_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(106),
	TestSignalName => "MCMIREADDATA(106)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(106),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(106),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(106),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(106),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(106),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA107_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA107_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(107),
	TestSignalName => "MCMIREADDATA(107)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(107),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(107),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(107),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(107),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(107),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA108_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA108_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(108),
	TestSignalName => "MCMIREADDATA(108)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(108),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(108),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(108),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(108),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(108),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA109_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA109_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(109),
	TestSignalName => "MCMIREADDATA(109)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(109),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(109),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(109),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(109),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(109),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA110_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA110_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(110),
	TestSignalName => "MCMIREADDATA(110)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(110),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(110),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(110),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(110),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(110),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA111_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA111_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(111),
	TestSignalName => "MCMIREADDATA(111)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(111),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(111),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(111),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(111),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(111),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA112_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA112_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(112),
	TestSignalName => "MCMIREADDATA(112)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(112),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(112),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(112),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(112),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(112),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA113_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA113_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(113),
	TestSignalName => "MCMIREADDATA(113)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(113),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(113),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(113),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(113),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(113),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA114_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA114_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(114),
	TestSignalName => "MCMIREADDATA(114)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(114),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(114),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(114),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(114),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(114),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA115_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA115_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(115),
	TestSignalName => "MCMIREADDATA(115)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(115),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(115),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(115),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(115),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(115),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA116_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA116_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(116),
	TestSignalName => "MCMIREADDATA(116)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(116),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(116),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(116),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(116),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(116),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA117_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA117_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(117),
	TestSignalName => "MCMIREADDATA(117)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(117),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(117),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(117),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(117),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(117),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA118_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA118_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(118),
	TestSignalName => "MCMIREADDATA(118)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(118),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(118),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(118),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(118),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(118),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA119_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA119_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(119),
	TestSignalName => "MCMIREADDATA(119)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(119),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(119),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(119),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(119),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(119),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA120_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA120_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(120),
	TestSignalName => "MCMIREADDATA(120)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(120),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(120),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(120),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(120),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(120),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA121_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA121_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(121),
	TestSignalName => "MCMIREADDATA(121)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(121),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(121),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(121),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(121),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(121),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA122_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA122_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(122),
	TestSignalName => "MCMIREADDATA(122)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(122),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(122),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(122),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(122),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(122),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA123_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA123_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(123),
	TestSignalName => "MCMIREADDATA(123)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(123),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(123),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(123),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(123),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(123),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA124_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA124_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(124),
	TestSignalName => "MCMIREADDATA(124)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(124),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(124),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(124),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(124),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(124),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA125_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA125_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(125),
	TestSignalName => "MCMIREADDATA(125)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(125),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(125),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(125),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(125),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(125),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA126_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA126_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(126),
	TestSignalName => "MCMIREADDATA(126)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(126),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(126),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(126),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(126),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(126),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation => Tviol_MCMIREADDATA127_CPMMCCLK_posedge,
	TimingData => Tmkr_MCMIREADDATA127_CPMMCCLK_posedge,
	TestSignal => MCMIREADDATA_dly(127),
	TestSignalName => "MCMIREADDATA(127)",
	TestDelay => tisd_MCMIREADDATA_CPMMCCLK(127),
	RefSignal => CPMMCCLK_dly,
	RefSignalName => "CPMMCCLK",
	RefDelay => ticd_CPMMCCLK,
	SetupHigh => tsetup_MCMIREADDATA_CPMMCCLK_posedge_posedge(127),
	SetupLow => tsetup_MCMIREADDATA_CPMMCCLK_negedge_posedge(127),
	HoldLow => thold_MCMIREADDATA_CPMMCCLK_posedge_posedge(127),
	HoldHigh => thold_MCMIREADDATA_CPMMCCLK_negedge_posedge(127),
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_MCMIREADDATAERR_CPMMCCLK_posedge,
	TimingData     => Tmkr_MCMIREADDATAERR_CPMMCCLK_posedge,
	TestSignal     => MCMIREADDATAERR,
	TestSignalName => "MCMIREADDATAERR",
	TestDelay      => 0 ps,
	RefSignal => CPMMCCLK_dly,
	RefSignalName  => "CPMMCCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_MCMIREADDATAERR_CPMMCCLK_posedge_posedge,
	SetupLow       => tsetup_MCMIREADDATAERR_CPMMCCLK_negedge_posedge,
	HoldLow        => thold_MCMIREADDATAERR_CPMMCCLK_posedge_posedge,
	HoldHigh       => thold_MCMIREADDATAERR_CPMMCCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_MCMIREADDATAVALID_CPMMCCLK_posedge,
	TimingData     => Tmkr_MCMIREADDATAVALID_CPMMCCLK_posedge,
	TestSignal     => MCMIREADDATAVALID,
	TestSignalName => "MCMIREADDATAVALID",
	TestDelay      => 0 ps,
	RefSignal => CPMMCCLK_dly,
	RefSignalName  => "CPMMCCLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_MCMIREADDATAVALID_CPMMCCLK_posedge_posedge,
	SetupLow       => tsetup_MCMIREADDATAVALID_CPMMCCLK_negedge_posedge,
	HoldLow        => thold_MCMIREADDATAVALID_CPMMCCLK_posedge_posedge,
	HoldHigh       => thold_MCMIREADDATAVALID_CPMMCCLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_TRCC440TRACEDISABLE_CPMC440CLK_posedge,
	TimingData     => Tmkr_TRCC440TRACEDISABLE_CPMC440CLK_posedge,
	TestSignal     => TRCC440TRACEDISABLE,
	TestSignalName => "TRCC440TRACEDISABLE",
	TestDelay      => 0 ps,
	RefSignal => CPMC440CLK_dly,
	RefSignalName  => "CPMC440CLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_TRCC440TRACEDISABLE_CPMC440CLK_posedge_posedge,
	SetupLow       => tsetup_TRCC440TRACEDISABLE_CPMC440CLK_negedge_posedge,
	HoldLow        => thold_TRCC440TRACEDISABLE_CPMC440CLK_posedge_posedge,
	HoldHigh       => thold_TRCC440TRACEDISABLE_CPMC440CLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
	VitalSetupHoldCheck
	(
	Violation      => Tviol_TRCC440TRIGGEREVENTIN_CPMC440CLK_posedge,
	TimingData     => Tmkr_TRCC440TRIGGEREVENTIN_CPMC440CLK_posedge,
	TestSignal     => TRCC440TRIGGEREVENTIN,
	TestSignalName => "TRCC440TRIGGEREVENTIN",
	TestDelay      => 0 ps,
	RefSignal => CPMC440CLK_dly,
	RefSignalName  => "CPMC440CLK",
	RefDelay       => 0 ps,
	SetupHigh      => tsetup_TRCC440TRIGGEREVENTIN_CPMC440CLK_posedge_posedge,
	SetupLow       => tsetup_TRCC440TRIGGEREVENTIN_CPMC440CLK_negedge_posedge,
	HoldLow        => thold_TRCC440TRIGGEREVENTIN_CPMC440CLK_posedge_posedge,
	HoldHigh       => thold_TRCC440TRIGGEREVENTIN_CPMC440CLK_negedge_posedge,
	CheckEnabled   => TRUE,
	RefTransition  => 'R',
	HeaderMsg      => InstancePath & "/X_PPC440",
	Xon            => Xon,
	MsgOn          => MsgOn,
	MsgSeverity    => WARNING
	);
     end if;
	VitalPathDelay01
	(
	OutSignal     => DMA0LLRSTENGINEACK,
	GlitchData    => DMA0LLRSTENGINEACK_GlitchData,
	OutSignalName => "DMA0LLRSTENGINEACK",
	OutTemp       => DMA0LLRSTENGINEACK_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLRSTENGINEACK,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLRSTENGINEACK, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLRXDSTRDYN,
	GlitchData    => DMA0LLRXDSTRDYN_GlitchData,
	OutSignalName => "DMA0LLRXDSTRDYN",
	OutTemp       => DMA0LLRXDSTRDYN_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLRXDSTRDYN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLRXDSTRDYN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(0),
	GlitchData    => DMA0LLTXD0_GlitchData,
	OutSignalName => "DMA0LLTXD(0)",
	OutTemp       => DMA0LLTXD_OUT(0),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(0),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(1),
	GlitchData    => DMA0LLTXD1_GlitchData,
	OutSignalName => "DMA0LLTXD(1)",
	OutTemp       => DMA0LLTXD_OUT(1),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(1),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(2),
	GlitchData    => DMA0LLTXD2_GlitchData,
	OutSignalName => "DMA0LLTXD(2)",
	OutTemp       => DMA0LLTXD_OUT(2),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(2),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(3),
	GlitchData    => DMA0LLTXD3_GlitchData,
	OutSignalName => "DMA0LLTXD(3)",
	OutTemp       => DMA0LLTXD_OUT(3),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(3),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(4),
	GlitchData    => DMA0LLTXD4_GlitchData,
	OutSignalName => "DMA0LLTXD(4)",
	OutTemp       => DMA0LLTXD_OUT(4),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(4),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(5),
	GlitchData    => DMA0LLTXD5_GlitchData,
	OutSignalName => "DMA0LLTXD(5)",
	OutTemp       => DMA0LLTXD_OUT(5),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(5),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(6),
	GlitchData    => DMA0LLTXD6_GlitchData,
	OutSignalName => "DMA0LLTXD(6)",
	OutTemp       => DMA0LLTXD_OUT(6),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(6),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(7),
	GlitchData    => DMA0LLTXD7_GlitchData,
	OutSignalName => "DMA0LLTXD(7)",
	OutTemp       => DMA0LLTXD_OUT(7),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(7),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(8),
	GlitchData    => DMA0LLTXD8_GlitchData,
	OutSignalName => "DMA0LLTXD(8)",
	OutTemp       => DMA0LLTXD_OUT(8),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(8),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(9),
	GlitchData    => DMA0LLTXD9_GlitchData,
	OutSignalName => "DMA0LLTXD(9)",
	OutTemp       => DMA0LLTXD_OUT(9),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(9),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(10),
	GlitchData    => DMA0LLTXD10_GlitchData,
	OutSignalName => "DMA0LLTXD(10)",
	OutTemp       => DMA0LLTXD_OUT(10),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(10),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(11),
	GlitchData    => DMA0LLTXD11_GlitchData,
	OutSignalName => "DMA0LLTXD(11)",
	OutTemp       => DMA0LLTXD_OUT(11),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(11),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(12),
	GlitchData    => DMA0LLTXD12_GlitchData,
	OutSignalName => "DMA0LLTXD(12)",
	OutTemp       => DMA0LLTXD_OUT(12),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(12),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(13),
	GlitchData    => DMA0LLTXD13_GlitchData,
	OutSignalName => "DMA0LLTXD(13)",
	OutTemp       => DMA0LLTXD_OUT(13),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(13),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(14),
	GlitchData    => DMA0LLTXD14_GlitchData,
	OutSignalName => "DMA0LLTXD(14)",
	OutTemp       => DMA0LLTXD_OUT(14),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(14),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(15),
	GlitchData    => DMA0LLTXD15_GlitchData,
	OutSignalName => "DMA0LLTXD(15)",
	OutTemp       => DMA0LLTXD_OUT(15),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(15),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(16),
	GlitchData    => DMA0LLTXD16_GlitchData,
	OutSignalName => "DMA0LLTXD(16)",
	OutTemp       => DMA0LLTXD_OUT(16),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(16),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(17),
	GlitchData    => DMA0LLTXD17_GlitchData,
	OutSignalName => "DMA0LLTXD(17)",
	OutTemp       => DMA0LLTXD_OUT(17),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(17),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(18),
	GlitchData    => DMA0LLTXD18_GlitchData,
	OutSignalName => "DMA0LLTXD(18)",
	OutTemp       => DMA0LLTXD_OUT(18),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(18),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(19),
	GlitchData    => DMA0LLTXD19_GlitchData,
	OutSignalName => "DMA0LLTXD(19)",
	OutTemp       => DMA0LLTXD_OUT(19),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(19),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(20),
	GlitchData    => DMA0LLTXD20_GlitchData,
	OutSignalName => "DMA0LLTXD(20)",
	OutTemp       => DMA0LLTXD_OUT(20),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(20),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(21),
	GlitchData    => DMA0LLTXD21_GlitchData,
	OutSignalName => "DMA0LLTXD(21)",
	OutTemp       => DMA0LLTXD_OUT(21),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(21),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(22),
	GlitchData    => DMA0LLTXD22_GlitchData,
	OutSignalName => "DMA0LLTXD(22)",
	OutTemp       => DMA0LLTXD_OUT(22),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(22),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(23),
	GlitchData    => DMA0LLTXD23_GlitchData,
	OutSignalName => "DMA0LLTXD(23)",
	OutTemp       => DMA0LLTXD_OUT(23),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(23),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(24),
	GlitchData    => DMA0LLTXD24_GlitchData,
	OutSignalName => "DMA0LLTXD(24)",
	OutTemp       => DMA0LLTXD_OUT(24),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(24),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(25),
	GlitchData    => DMA0LLTXD25_GlitchData,
	OutSignalName => "DMA0LLTXD(25)",
	OutTemp       => DMA0LLTXD_OUT(25),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(25),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(26),
	GlitchData    => DMA0LLTXD26_GlitchData,
	OutSignalName => "DMA0LLTXD(26)",
	OutTemp       => DMA0LLTXD_OUT(26),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(26),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(27),
	GlitchData    => DMA0LLTXD27_GlitchData,
	OutSignalName => "DMA0LLTXD(27)",
	OutTemp       => DMA0LLTXD_OUT(27),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(27),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(28),
	GlitchData    => DMA0LLTXD28_GlitchData,
	OutSignalName => "DMA0LLTXD(28)",
	OutTemp       => DMA0LLTXD_OUT(28),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(28),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(29),
	GlitchData    => DMA0LLTXD29_GlitchData,
	OutSignalName => "DMA0LLTXD(29)",
	OutTemp       => DMA0LLTXD_OUT(29),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(29),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(30),
	GlitchData    => DMA0LLTXD30_GlitchData,
	OutSignalName => "DMA0LLTXD(30)",
	OutTemp       => DMA0LLTXD_OUT(30),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(30),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXD(31),
	GlitchData    => DMA0LLTXD31_GlitchData,
	OutSignalName => "DMA0LLTXD(31)",
	OutTemp       => DMA0LLTXD_OUT(31),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXD(31),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXD(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXEOFN,
	GlitchData    => DMA0LLTXEOFN_GlitchData,
	OutSignalName => "DMA0LLTXEOFN",
	OutTemp       => DMA0LLTXEOFN_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXEOFN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXEOFN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXEOPN,
	GlitchData    => DMA0LLTXEOPN_GlitchData,
	OutSignalName => "DMA0LLTXEOPN",
	OutTemp       => DMA0LLTXEOPN_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXEOPN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXEOPN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXREM(0),
	GlitchData    => DMA0LLTXREM0_GlitchData,
	OutSignalName => "DMA0LLTXREM(0)",
	OutTemp       => DMA0LLTXREM_OUT(0),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXREM(0),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXREM(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXREM(1),
	GlitchData    => DMA0LLTXREM1_GlitchData,
	OutSignalName => "DMA0LLTXREM(1)",
	OutTemp       => DMA0LLTXREM_OUT(1),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXREM(1),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXREM(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXREM(2),
	GlitchData    => DMA0LLTXREM2_GlitchData,
	OutSignalName => "DMA0LLTXREM(2)",
	OutTemp       => DMA0LLTXREM_OUT(2),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXREM(2),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXREM(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXREM(3),
	GlitchData    => DMA0LLTXREM3_GlitchData,
	OutSignalName => "DMA0LLTXREM(3)",
	OutTemp       => DMA0LLTXREM_OUT(3),
	Paths       => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXREM(3),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXREM(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXSOFN,
	GlitchData    => DMA0LLTXSOFN_GlitchData,
	OutSignalName => "DMA0LLTXSOFN",
	OutTemp       => DMA0LLTXSOFN_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXSOFN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXSOFN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXSOPN,
	GlitchData    => DMA0LLTXSOPN_GlitchData,
	OutSignalName => "DMA0LLTXSOPN",
	OutTemp       => DMA0LLTXSOPN_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXSOPN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXSOPN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0LLTXSRCRDYN,
	GlitchData    => DMA0LLTXSRCRDYN_GlitchData,
	OutSignalName => "DMA0LLTXSRCRDYN",
	OutTemp       => DMA0LLTXSRCRDYN_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0LLTXSRCRDYN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0LLTXSRCRDYN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0RXIRQ,
	GlitchData    => DMA0RXIRQ_GlitchData,
	OutSignalName => "DMA0RXIRQ",
	OutTemp       => DMA0RXIRQ_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0RXIRQ,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0RXIRQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA0TXIRQ,
	GlitchData    => DMA0TXIRQ_GlitchData,
	OutSignalName => "DMA0TXIRQ",
	OutTemp       => DMA0TXIRQ_OUT,
	Paths         => (0 => (CPMDMA0LLCLK_dly'last_event, tpd_CPMDMA0LLCLK_DMA0TXIRQ,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA0LLCLK_DMA0TXIRQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLRSTENGINEACK,
	GlitchData    => DMA1LLRSTENGINEACK_GlitchData,
	OutSignalName => "DMA1LLRSTENGINEACK",
	OutTemp       => DMA1LLRSTENGINEACK_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLRSTENGINEACK,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLRSTENGINEACK, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLRXDSTRDYN,
	GlitchData    => DMA1LLRXDSTRDYN_GlitchData,
	OutSignalName => "DMA1LLRXDSTRDYN",
	OutTemp       => DMA1LLRXDSTRDYN_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLRXDSTRDYN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLRXDSTRDYN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(0),
	GlitchData    => DMA1LLTXD0_GlitchData,
	OutSignalName => "DMA1LLTXD(0)",
	OutTemp       => DMA1LLTXD_OUT(0),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(0),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(1),
	GlitchData    => DMA1LLTXD1_GlitchData,
	OutSignalName => "DMA1LLTXD(1)",
	OutTemp       => DMA1LLTXD_OUT(1),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(1),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(2),
	GlitchData    => DMA1LLTXD2_GlitchData,
	OutSignalName => "DMA1LLTXD(2)",
	OutTemp       => DMA1LLTXD_OUT(2),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(2),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(3),
	GlitchData    => DMA1LLTXD3_GlitchData,
	OutSignalName => "DMA1LLTXD(3)",
	OutTemp       => DMA1LLTXD_OUT(3),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(3),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(4),
	GlitchData    => DMA1LLTXD4_GlitchData,
	OutSignalName => "DMA1LLTXD(4)",
	OutTemp       => DMA1LLTXD_OUT(4),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(4),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(5),
	GlitchData    => DMA1LLTXD5_GlitchData,
	OutSignalName => "DMA1LLTXD(5)",
	OutTemp       => DMA1LLTXD_OUT(5),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(5),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(6),
	GlitchData    => DMA1LLTXD6_GlitchData,
	OutSignalName => "DMA1LLTXD(6)",
	OutTemp       => DMA1LLTXD_OUT(6),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(6),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(7),
	GlitchData    => DMA1LLTXD7_GlitchData,
	OutSignalName => "DMA1LLTXD(7)",
	OutTemp       => DMA1LLTXD_OUT(7),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(7),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(8),
	GlitchData    => DMA1LLTXD8_GlitchData,
	OutSignalName => "DMA1LLTXD(8)",
	OutTemp       => DMA1LLTXD_OUT(8),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(8),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(9),
	GlitchData    => DMA1LLTXD9_GlitchData,
	OutSignalName => "DMA1LLTXD(9)",
	OutTemp       => DMA1LLTXD_OUT(9),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(9),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(10),
	GlitchData    => DMA1LLTXD10_GlitchData,
	OutSignalName => "DMA1LLTXD(10)",
	OutTemp       => DMA1LLTXD_OUT(10),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(10),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(11),
	GlitchData    => DMA1LLTXD11_GlitchData,
	OutSignalName => "DMA1LLTXD(11)",
	OutTemp       => DMA1LLTXD_OUT(11),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(11),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(12),
	GlitchData    => DMA1LLTXD12_GlitchData,
	OutSignalName => "DMA1LLTXD(12)",
	OutTemp       => DMA1LLTXD_OUT(12),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(12),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(13),
	GlitchData    => DMA1LLTXD13_GlitchData,
	OutSignalName => "DMA1LLTXD(13)",
	OutTemp       => DMA1LLTXD_OUT(13),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(13),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(14),
	GlitchData    => DMA1LLTXD14_GlitchData,
	OutSignalName => "DMA1LLTXD(14)",
	OutTemp       => DMA1LLTXD_OUT(14),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(14),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(15),
	GlitchData    => DMA1LLTXD15_GlitchData,
	OutSignalName => "DMA1LLTXD(15)",
	OutTemp       => DMA1LLTXD_OUT(15),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(15),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(16),
	GlitchData    => DMA1LLTXD16_GlitchData,
	OutSignalName => "DMA1LLTXD(16)",
	OutTemp       => DMA1LLTXD_OUT(16),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(16),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(17),
	GlitchData    => DMA1LLTXD17_GlitchData,
	OutSignalName => "DMA1LLTXD(17)",
	OutTemp       => DMA1LLTXD_OUT(17),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(17),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(18),
	GlitchData    => DMA1LLTXD18_GlitchData,
	OutSignalName => "DMA1LLTXD(18)",
	OutTemp       => DMA1LLTXD_OUT(18),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(18),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(19),
	GlitchData    => DMA1LLTXD19_GlitchData,
	OutSignalName => "DMA1LLTXD(19)",
	OutTemp       => DMA1LLTXD_OUT(19),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(19),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(20),
	GlitchData    => DMA1LLTXD20_GlitchData,
	OutSignalName => "DMA1LLTXD(20)",
	OutTemp       => DMA1LLTXD_OUT(20),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(20),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(21),
	GlitchData    => DMA1LLTXD21_GlitchData,
	OutSignalName => "DMA1LLTXD(21)",
	OutTemp       => DMA1LLTXD_OUT(21),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(21),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(22),
	GlitchData    => DMA1LLTXD22_GlitchData,
	OutSignalName => "DMA1LLTXD(22)",
	OutTemp       => DMA1LLTXD_OUT(22),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(22),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(23),
	GlitchData    => DMA1LLTXD23_GlitchData,
	OutSignalName => "DMA1LLTXD(23)",
	OutTemp       => DMA1LLTXD_OUT(23),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(23),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(24),
	GlitchData    => DMA1LLTXD24_GlitchData,
	OutSignalName => "DMA1LLTXD(24)",
	OutTemp       => DMA1LLTXD_OUT(24),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(24),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(25),
	GlitchData    => DMA1LLTXD25_GlitchData,
	OutSignalName => "DMA1LLTXD(25)",
	OutTemp       => DMA1LLTXD_OUT(25),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(25),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(26),
	GlitchData    => DMA1LLTXD26_GlitchData,
	OutSignalName => "DMA1LLTXD(26)",
	OutTemp       => DMA1LLTXD_OUT(26),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(26),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(27),
	GlitchData    => DMA1LLTXD27_GlitchData,
	OutSignalName => "DMA1LLTXD(27)",
	OutTemp       => DMA1LLTXD_OUT(27),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(27),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(28),
	GlitchData    => DMA1LLTXD28_GlitchData,
	OutSignalName => "DMA1LLTXD(28)",
	OutTemp       => DMA1LLTXD_OUT(28),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(28),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(29),
	GlitchData    => DMA1LLTXD29_GlitchData,
	OutSignalName => "DMA1LLTXD(29)",
	OutTemp       => DMA1LLTXD_OUT(29),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(29),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(30),
	GlitchData    => DMA1LLTXD30_GlitchData,
	OutSignalName => "DMA1LLTXD(30)",
	OutTemp       => DMA1LLTXD_OUT(30),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(30),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXD(31),
	GlitchData    => DMA1LLTXD31_GlitchData,
	OutSignalName => "DMA1LLTXD(31)",
	OutTemp       => DMA1LLTXD_OUT(31),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXD(31),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXD(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXEOFN,
	GlitchData    => DMA1LLTXEOFN_GlitchData,
	OutSignalName => "DMA1LLTXEOFN",
	OutTemp       => DMA1LLTXEOFN_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXEOFN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXEOFN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXEOPN,
	GlitchData    => DMA1LLTXEOPN_GlitchData,
	OutSignalName => "DMA1LLTXEOPN",
	OutTemp       => DMA1LLTXEOPN_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXEOPN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXEOPN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXREM(0),
	GlitchData    => DMA1LLTXREM0_GlitchData,
	OutSignalName => "DMA1LLTXREM(0)",
	OutTemp       => DMA1LLTXREM_OUT(0),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXREM(0),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXREM(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXREM(1),
	GlitchData    => DMA1LLTXREM1_GlitchData,
	OutSignalName => "DMA1LLTXREM(1)",
	OutTemp       => DMA1LLTXREM_OUT(1),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXREM(1),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXREM(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXREM(2),
	GlitchData    => DMA1LLTXREM2_GlitchData,
	OutSignalName => "DMA1LLTXREM(2)",
	OutTemp       => DMA1LLTXREM_OUT(2),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXREM(2),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXREM(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXREM(3),
	GlitchData    => DMA1LLTXREM3_GlitchData,
	OutSignalName => "DMA1LLTXREM(3)",
	OutTemp       => DMA1LLTXREM_OUT(3),
	Paths       => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXREM(3),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXREM(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXSOFN,
	GlitchData    => DMA1LLTXSOFN_GlitchData,
	OutSignalName => "DMA1LLTXSOFN",
	OutTemp       => DMA1LLTXSOFN_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXSOFN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXSOFN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXSOPN,
	GlitchData    => DMA1LLTXSOPN_GlitchData,
	OutSignalName => "DMA1LLTXSOPN",
	OutTemp       => DMA1LLTXSOPN_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXSOPN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXSOPN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1LLTXSRCRDYN,
	GlitchData    => DMA1LLTXSRCRDYN_GlitchData,
	OutSignalName => "DMA1LLTXSRCRDYN",
	OutTemp       => DMA1LLTXSRCRDYN_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1LLTXSRCRDYN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1LLTXSRCRDYN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1RXIRQ,
	GlitchData    => DMA1RXIRQ_GlitchData,
	OutSignalName => "DMA1RXIRQ",
	OutTemp       => DMA1RXIRQ_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1RXIRQ,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1RXIRQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA1TXIRQ,
	GlitchData    => DMA1TXIRQ_GlitchData,
	OutSignalName => "DMA1TXIRQ",
	OutTemp       => DMA1TXIRQ_OUT,
	Paths         => (0 => (CPMDMA1LLCLK_dly'last_event, tpd_CPMDMA1LLCLK_DMA1TXIRQ,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA1LLCLK_DMA1TXIRQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLRSTENGINEACK,
	GlitchData    => DMA2LLRSTENGINEACK_GlitchData,
	OutSignalName => "DMA2LLRSTENGINEACK",
	OutTemp       => DMA2LLRSTENGINEACK_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLRSTENGINEACK,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLRSTENGINEACK, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLRXDSTRDYN,
	GlitchData    => DMA2LLRXDSTRDYN_GlitchData,
	OutSignalName => "DMA2LLRXDSTRDYN",
	OutTemp       => DMA2LLRXDSTRDYN_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLRXDSTRDYN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLRXDSTRDYN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(0),
	GlitchData    => DMA2LLTXD0_GlitchData,
	OutSignalName => "DMA2LLTXD(0)",
	OutTemp       => DMA2LLTXD_OUT(0),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(0),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(1),
	GlitchData    => DMA2LLTXD1_GlitchData,
	OutSignalName => "DMA2LLTXD(1)",
	OutTemp       => DMA2LLTXD_OUT(1),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(1),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(2),
	GlitchData    => DMA2LLTXD2_GlitchData,
	OutSignalName => "DMA2LLTXD(2)",
	OutTemp       => DMA2LLTXD_OUT(2),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(2),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(3),
	GlitchData    => DMA2LLTXD3_GlitchData,
	OutSignalName => "DMA2LLTXD(3)",
	OutTemp       => DMA2LLTXD_OUT(3),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(3),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(4),
	GlitchData    => DMA2LLTXD4_GlitchData,
	OutSignalName => "DMA2LLTXD(4)",
	OutTemp       => DMA2LLTXD_OUT(4),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(4),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(5),
	GlitchData    => DMA2LLTXD5_GlitchData,
	OutSignalName => "DMA2LLTXD(5)",
	OutTemp       => DMA2LLTXD_OUT(5),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(5),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(6),
	GlitchData    => DMA2LLTXD6_GlitchData,
	OutSignalName => "DMA2LLTXD(6)",
	OutTemp       => DMA2LLTXD_OUT(6),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(6),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(7),
	GlitchData    => DMA2LLTXD7_GlitchData,
	OutSignalName => "DMA2LLTXD(7)",
	OutTemp       => DMA2LLTXD_OUT(7),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(7),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(8),
	GlitchData    => DMA2LLTXD8_GlitchData,
	OutSignalName => "DMA2LLTXD(8)",
	OutTemp       => DMA2LLTXD_OUT(8),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(8),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(9),
	GlitchData    => DMA2LLTXD9_GlitchData,
	OutSignalName => "DMA2LLTXD(9)",
	OutTemp       => DMA2LLTXD_OUT(9),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(9),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(10),
	GlitchData    => DMA2LLTXD10_GlitchData,
	OutSignalName => "DMA2LLTXD(10)",
	OutTemp       => DMA2LLTXD_OUT(10),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(10),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(11),
	GlitchData    => DMA2LLTXD11_GlitchData,
	OutSignalName => "DMA2LLTXD(11)",
	OutTemp       => DMA2LLTXD_OUT(11),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(11),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(12),
	GlitchData    => DMA2LLTXD12_GlitchData,
	OutSignalName => "DMA2LLTXD(12)",
	OutTemp       => DMA2LLTXD_OUT(12),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(12),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(13),
	GlitchData    => DMA2LLTXD13_GlitchData,
	OutSignalName => "DMA2LLTXD(13)",
	OutTemp       => DMA2LLTXD_OUT(13),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(13),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(14),
	GlitchData    => DMA2LLTXD14_GlitchData,
	OutSignalName => "DMA2LLTXD(14)",
	OutTemp       => DMA2LLTXD_OUT(14),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(14),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(15),
	GlitchData    => DMA2LLTXD15_GlitchData,
	OutSignalName => "DMA2LLTXD(15)",
	OutTemp       => DMA2LLTXD_OUT(15),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(15),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(16),
	GlitchData    => DMA2LLTXD16_GlitchData,
	OutSignalName => "DMA2LLTXD(16)",
	OutTemp       => DMA2LLTXD_OUT(16),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(16),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(17),
	GlitchData    => DMA2LLTXD17_GlitchData,
	OutSignalName => "DMA2LLTXD(17)",
	OutTemp       => DMA2LLTXD_OUT(17),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(17),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(18),
	GlitchData    => DMA2LLTXD18_GlitchData,
	OutSignalName => "DMA2LLTXD(18)",
	OutTemp       => DMA2LLTXD_OUT(18),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(18),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(19),
	GlitchData    => DMA2LLTXD19_GlitchData,
	OutSignalName => "DMA2LLTXD(19)",
	OutTemp       => DMA2LLTXD_OUT(19),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(19),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(20),
	GlitchData    => DMA2LLTXD20_GlitchData,
	OutSignalName => "DMA2LLTXD(20)",
	OutTemp       => DMA2LLTXD_OUT(20),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(20),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(21),
	GlitchData    => DMA2LLTXD21_GlitchData,
	OutSignalName => "DMA2LLTXD(21)",
	OutTemp       => DMA2LLTXD_OUT(21),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(21),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(22),
	GlitchData    => DMA2LLTXD22_GlitchData,
	OutSignalName => "DMA2LLTXD(22)",
	OutTemp       => DMA2LLTXD_OUT(22),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(22),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(23),
	GlitchData    => DMA2LLTXD23_GlitchData,
	OutSignalName => "DMA2LLTXD(23)",
	OutTemp       => DMA2LLTXD_OUT(23),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(23),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(24),
	GlitchData    => DMA2LLTXD24_GlitchData,
	OutSignalName => "DMA2LLTXD(24)",
	OutTemp       => DMA2LLTXD_OUT(24),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(24),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(25),
	GlitchData    => DMA2LLTXD25_GlitchData,
	OutSignalName => "DMA2LLTXD(25)",
	OutTemp       => DMA2LLTXD_OUT(25),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(25),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(26),
	GlitchData    => DMA2LLTXD26_GlitchData,
	OutSignalName => "DMA2LLTXD(26)",
	OutTemp       => DMA2LLTXD_OUT(26),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(26),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(27),
	GlitchData    => DMA2LLTXD27_GlitchData,
	OutSignalName => "DMA2LLTXD(27)",
	OutTemp       => DMA2LLTXD_OUT(27),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(27),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(28),
	GlitchData    => DMA2LLTXD28_GlitchData,
	OutSignalName => "DMA2LLTXD(28)",
	OutTemp       => DMA2LLTXD_OUT(28),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(28),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(29),
	GlitchData    => DMA2LLTXD29_GlitchData,
	OutSignalName => "DMA2LLTXD(29)",
	OutTemp       => DMA2LLTXD_OUT(29),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(29),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(30),
	GlitchData    => DMA2LLTXD30_GlitchData,
	OutSignalName => "DMA2LLTXD(30)",
	OutTemp       => DMA2LLTXD_OUT(30),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(30),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXD(31),
	GlitchData    => DMA2LLTXD31_GlitchData,
	OutSignalName => "DMA2LLTXD(31)",
	OutTemp       => DMA2LLTXD_OUT(31),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXD(31),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXD(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXEOFN,
	GlitchData    => DMA2LLTXEOFN_GlitchData,
	OutSignalName => "DMA2LLTXEOFN",
	OutTemp       => DMA2LLTXEOFN_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXEOFN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXEOFN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXEOPN,
	GlitchData    => DMA2LLTXEOPN_GlitchData,
	OutSignalName => "DMA2LLTXEOPN",
	OutTemp       => DMA2LLTXEOPN_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXEOPN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXEOPN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXREM(0),
	GlitchData    => DMA2LLTXREM0_GlitchData,
	OutSignalName => "DMA2LLTXREM(0)",
	OutTemp       => DMA2LLTXREM_OUT(0),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXREM(0),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXREM(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXREM(1),
	GlitchData    => DMA2LLTXREM1_GlitchData,
	OutSignalName => "DMA2LLTXREM(1)",
	OutTemp       => DMA2LLTXREM_OUT(1),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXREM(1),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXREM(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXREM(2),
	GlitchData    => DMA2LLTXREM2_GlitchData,
	OutSignalName => "DMA2LLTXREM(2)",
	OutTemp       => DMA2LLTXREM_OUT(2),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXREM(2),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXREM(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXREM(3),
	GlitchData    => DMA2LLTXREM3_GlitchData,
	OutSignalName => "DMA2LLTXREM(3)",
	OutTemp       => DMA2LLTXREM_OUT(3),
	Paths       => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXREM(3),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXREM(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXSOFN,
	GlitchData    => DMA2LLTXSOFN_GlitchData,
	OutSignalName => "DMA2LLTXSOFN",
	OutTemp       => DMA2LLTXSOFN_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXSOFN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXSOFN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXSOPN,
	GlitchData    => DMA2LLTXSOPN_GlitchData,
	OutSignalName => "DMA2LLTXSOPN",
	OutTemp       => DMA2LLTXSOPN_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXSOPN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXSOPN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2LLTXSRCRDYN,
	GlitchData    => DMA2LLTXSRCRDYN_GlitchData,
	OutSignalName => "DMA2LLTXSRCRDYN",
	OutTemp       => DMA2LLTXSRCRDYN_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2LLTXSRCRDYN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2LLTXSRCRDYN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2RXIRQ,
	GlitchData    => DMA2RXIRQ_GlitchData,
	OutSignalName => "DMA2RXIRQ",
	OutTemp       => DMA2RXIRQ_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2RXIRQ,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2RXIRQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA2TXIRQ,
	GlitchData    => DMA2TXIRQ_GlitchData,
	OutSignalName => "DMA2TXIRQ",
	OutTemp       => DMA2TXIRQ_OUT,
	Paths         => (0 => (CPMDMA2LLCLK_dly'last_event, tpd_CPMDMA2LLCLK_DMA2TXIRQ,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA2LLCLK_DMA2TXIRQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLRSTENGINEACK,
	GlitchData    => DMA3LLRSTENGINEACK_GlitchData,
	OutSignalName => "DMA3LLRSTENGINEACK",
	OutTemp       => DMA3LLRSTENGINEACK_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLRSTENGINEACK,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLRSTENGINEACK, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLRXDSTRDYN,
	GlitchData    => DMA3LLRXDSTRDYN_GlitchData,
	OutSignalName => "DMA3LLRXDSTRDYN",
	OutTemp       => DMA3LLRXDSTRDYN_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLRXDSTRDYN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLRXDSTRDYN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(0),
	GlitchData    => DMA3LLTXD0_GlitchData,
	OutSignalName => "DMA3LLTXD(0)",
	OutTemp       => DMA3LLTXD_OUT(0),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(0),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(1),
	GlitchData    => DMA3LLTXD1_GlitchData,
	OutSignalName => "DMA3LLTXD(1)",
	OutTemp       => DMA3LLTXD_OUT(1),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(1),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(2),
	GlitchData    => DMA3LLTXD2_GlitchData,
	OutSignalName => "DMA3LLTXD(2)",
	OutTemp       => DMA3LLTXD_OUT(2),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(2),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(3),
	GlitchData    => DMA3LLTXD3_GlitchData,
	OutSignalName => "DMA3LLTXD(3)",
	OutTemp       => DMA3LLTXD_OUT(3),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(3),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(4),
	GlitchData    => DMA3LLTXD4_GlitchData,
	OutSignalName => "DMA3LLTXD(4)",
	OutTemp       => DMA3LLTXD_OUT(4),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(4),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(5),
	GlitchData    => DMA3LLTXD5_GlitchData,
	OutSignalName => "DMA3LLTXD(5)",
	OutTemp       => DMA3LLTXD_OUT(5),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(5),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(6),
	GlitchData    => DMA3LLTXD6_GlitchData,
	OutSignalName => "DMA3LLTXD(6)",
	OutTemp       => DMA3LLTXD_OUT(6),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(6),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(7),
	GlitchData    => DMA3LLTXD7_GlitchData,
	OutSignalName => "DMA3LLTXD(7)",
	OutTemp       => DMA3LLTXD_OUT(7),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(7),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(8),
	GlitchData    => DMA3LLTXD8_GlitchData,
	OutSignalName => "DMA3LLTXD(8)",
	OutTemp       => DMA3LLTXD_OUT(8),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(8),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(9),
	GlitchData    => DMA3LLTXD9_GlitchData,
	OutSignalName => "DMA3LLTXD(9)",
	OutTemp       => DMA3LLTXD_OUT(9),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(9),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(10),
	GlitchData    => DMA3LLTXD10_GlitchData,
	OutSignalName => "DMA3LLTXD(10)",
	OutTemp       => DMA3LLTXD_OUT(10),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(10),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(11),
	GlitchData    => DMA3LLTXD11_GlitchData,
	OutSignalName => "DMA3LLTXD(11)",
	OutTemp       => DMA3LLTXD_OUT(11),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(11),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(12),
	GlitchData    => DMA3LLTXD12_GlitchData,
	OutSignalName => "DMA3LLTXD(12)",
	OutTemp       => DMA3LLTXD_OUT(12),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(12),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(13),
	GlitchData    => DMA3LLTXD13_GlitchData,
	OutSignalName => "DMA3LLTXD(13)",
	OutTemp       => DMA3LLTXD_OUT(13),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(13),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(14),
	GlitchData    => DMA3LLTXD14_GlitchData,
	OutSignalName => "DMA3LLTXD(14)",
	OutTemp       => DMA3LLTXD_OUT(14),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(14),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(15),
	GlitchData    => DMA3LLTXD15_GlitchData,
	OutSignalName => "DMA3LLTXD(15)",
	OutTemp       => DMA3LLTXD_OUT(15),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(15),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(16),
	GlitchData    => DMA3LLTXD16_GlitchData,
	OutSignalName => "DMA3LLTXD(16)",
	OutTemp       => DMA3LLTXD_OUT(16),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(16),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(17),
	GlitchData    => DMA3LLTXD17_GlitchData,
	OutSignalName => "DMA3LLTXD(17)",
	OutTemp       => DMA3LLTXD_OUT(17),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(17),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(18),
	GlitchData    => DMA3LLTXD18_GlitchData,
	OutSignalName => "DMA3LLTXD(18)",
	OutTemp       => DMA3LLTXD_OUT(18),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(18),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(19),
	GlitchData    => DMA3LLTXD19_GlitchData,
	OutSignalName => "DMA3LLTXD(19)",
	OutTemp       => DMA3LLTXD_OUT(19),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(19),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(20),
	GlitchData    => DMA3LLTXD20_GlitchData,
	OutSignalName => "DMA3LLTXD(20)",
	OutTemp       => DMA3LLTXD_OUT(20),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(20),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(21),
	GlitchData    => DMA3LLTXD21_GlitchData,
	OutSignalName => "DMA3LLTXD(21)",
	OutTemp       => DMA3LLTXD_OUT(21),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(21),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(22),
	GlitchData    => DMA3LLTXD22_GlitchData,
	OutSignalName => "DMA3LLTXD(22)",
	OutTemp       => DMA3LLTXD_OUT(22),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(22),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(23),
	GlitchData    => DMA3LLTXD23_GlitchData,
	OutSignalName => "DMA3LLTXD(23)",
	OutTemp       => DMA3LLTXD_OUT(23),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(23),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(24),
	GlitchData    => DMA3LLTXD24_GlitchData,
	OutSignalName => "DMA3LLTXD(24)",
	OutTemp       => DMA3LLTXD_OUT(24),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(24),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(25),
	GlitchData    => DMA3LLTXD25_GlitchData,
	OutSignalName => "DMA3LLTXD(25)",
	OutTemp       => DMA3LLTXD_OUT(25),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(25),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(26),
	GlitchData    => DMA3LLTXD26_GlitchData,
	OutSignalName => "DMA3LLTXD(26)",
	OutTemp       => DMA3LLTXD_OUT(26),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(26),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(27),
	GlitchData    => DMA3LLTXD27_GlitchData,
	OutSignalName => "DMA3LLTXD(27)",
	OutTemp       => DMA3LLTXD_OUT(27),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(27),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(28),
	GlitchData    => DMA3LLTXD28_GlitchData,
	OutSignalName => "DMA3LLTXD(28)",
	OutTemp       => DMA3LLTXD_OUT(28),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(28),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(29),
	GlitchData    => DMA3LLTXD29_GlitchData,
	OutSignalName => "DMA3LLTXD(29)",
	OutTemp       => DMA3LLTXD_OUT(29),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(29),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(30),
	GlitchData    => DMA3LLTXD30_GlitchData,
	OutSignalName => "DMA3LLTXD(30)",
	OutTemp       => DMA3LLTXD_OUT(30),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(30),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXD(31),
	GlitchData    => DMA3LLTXD31_GlitchData,
	OutSignalName => "DMA3LLTXD(31)",
	OutTemp       => DMA3LLTXD_OUT(31),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXD(31),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXD(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXEOFN,
	GlitchData    => DMA3LLTXEOFN_GlitchData,
	OutSignalName => "DMA3LLTXEOFN",
	OutTemp       => DMA3LLTXEOFN_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXEOFN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXEOFN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXEOPN,
	GlitchData    => DMA3LLTXEOPN_GlitchData,
	OutSignalName => "DMA3LLTXEOPN",
	OutTemp       => DMA3LLTXEOPN_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXEOPN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXEOPN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXREM(0),
	GlitchData    => DMA3LLTXREM0_GlitchData,
	OutSignalName => "DMA3LLTXREM(0)",
	OutTemp       => DMA3LLTXREM_OUT(0),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXREM(0),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXREM(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXREM(1),
	GlitchData    => DMA3LLTXREM1_GlitchData,
	OutSignalName => "DMA3LLTXREM(1)",
	OutTemp       => DMA3LLTXREM_OUT(1),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXREM(1),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXREM(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXREM(2),
	GlitchData    => DMA3LLTXREM2_GlitchData,
	OutSignalName => "DMA3LLTXREM(2)",
	OutTemp       => DMA3LLTXREM_OUT(2),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXREM(2),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXREM(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXREM(3),
	GlitchData    => DMA3LLTXREM3_GlitchData,
	OutSignalName => "DMA3LLTXREM(3)",
	OutTemp       => DMA3LLTXREM_OUT(3),
	Paths       => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXREM(3),TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXREM(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXSOFN,
	GlitchData    => DMA3LLTXSOFN_GlitchData,
	OutSignalName => "DMA3LLTXSOFN",
	OutTemp       => DMA3LLTXSOFN_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXSOFN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXSOFN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXSOPN,
	GlitchData    => DMA3LLTXSOPN_GlitchData,
	OutSignalName => "DMA3LLTXSOPN",
	OutTemp       => DMA3LLTXSOPN_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXSOPN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXSOPN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3LLTXSRCRDYN,
	GlitchData    => DMA3LLTXSRCRDYN_GlitchData,
	OutSignalName => "DMA3LLTXSRCRDYN",
	OutTemp       => DMA3LLTXSRCRDYN_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3LLTXSRCRDYN,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3LLTXSRCRDYN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3RXIRQ,
	GlitchData    => DMA3RXIRQ_GlitchData,
	OutSignalName => "DMA3RXIRQ",
	OutTemp       => DMA3RXIRQ_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3RXIRQ,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3RXIRQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => DMA3TXIRQ,
	GlitchData    => DMA3TXIRQ_GlitchData,
	OutSignalName => "DMA3TXIRQ",
	OutTemp       => DMA3TXIRQ_OUT,
	Paths         => (0 => (CPMDMA3LLCLK_dly'last_event, tpd_CPMDMA3LLCLK_DMA3TXIRQ,TRUE)),
	 DefaultDelay =>  tpd_CPMDMA3LLCLK_DMA3TXIRQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(0),
	GlitchData    => PPCDMDCRABUS0_GlitchData,
	OutSignalName => "PPCDMDCRABUS(0)",
	OutTemp       => PPCDMDCRABUS_OUT(0),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRABUS(0),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRABUS(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(1),
	GlitchData    => PPCDMDCRABUS1_GlitchData,
	OutSignalName => "PPCDMDCRABUS(1)",
	OutTemp       => PPCDMDCRABUS_OUT(1),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRABUS(1),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRABUS(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(2),
	GlitchData    => PPCDMDCRABUS2_GlitchData,
	OutSignalName => "PPCDMDCRABUS(2)",
	OutTemp       => PPCDMDCRABUS_OUT(2),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRABUS(2),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRABUS(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(3),
	GlitchData    => PPCDMDCRABUS3_GlitchData,
	OutSignalName => "PPCDMDCRABUS(3)",
	OutTemp       => PPCDMDCRABUS_OUT(3),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRABUS(3),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRABUS(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(4),
	GlitchData    => PPCDMDCRABUS4_GlitchData,
	OutSignalName => "PPCDMDCRABUS(4)",
	OutTemp       => PPCDMDCRABUS_OUT(4),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRABUS(4),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRABUS(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(5),
	GlitchData    => PPCDMDCRABUS5_GlitchData,
	OutSignalName => "PPCDMDCRABUS(5)",
	OutTemp       => PPCDMDCRABUS_OUT(5),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRABUS(5),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRABUS(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(6),
	GlitchData    => PPCDMDCRABUS6_GlitchData,
	OutSignalName => "PPCDMDCRABUS(6)",
	OutTemp       => PPCDMDCRABUS_OUT(6),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRABUS(6),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRABUS(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(7),
	GlitchData    => PPCDMDCRABUS7_GlitchData,
	OutSignalName => "PPCDMDCRABUS(7)",
	OutTemp       => PPCDMDCRABUS_OUT(7),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRABUS(7),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRABUS(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(8),
	GlitchData    => PPCDMDCRABUS8_GlitchData,
	OutSignalName => "PPCDMDCRABUS(8)",
	OutTemp       => PPCDMDCRABUS_OUT(8),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRABUS(8),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRABUS(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRABUS(9),
	GlitchData    => PPCDMDCRABUS9_GlitchData,
	OutSignalName => "PPCDMDCRABUS(9)",
	OutTemp       => PPCDMDCRABUS_OUT(9),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRABUS(9),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRABUS(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(0),
	GlitchData    => PPCDMDCRDBUSOUT0_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(0)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(0),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(0),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(1),
	GlitchData    => PPCDMDCRDBUSOUT1_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(1)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(1),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(1),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(2),
	GlitchData    => PPCDMDCRDBUSOUT2_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(2)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(2),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(2),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(3),
	GlitchData    => PPCDMDCRDBUSOUT3_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(3)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(3),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(3),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(4),
	GlitchData    => PPCDMDCRDBUSOUT4_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(4)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(4),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(4),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(5),
	GlitchData    => PPCDMDCRDBUSOUT5_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(5)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(5),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(5),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(6),
	GlitchData    => PPCDMDCRDBUSOUT6_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(6)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(6),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(6),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(7),
	GlitchData    => PPCDMDCRDBUSOUT7_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(7)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(7),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(7),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(8),
	GlitchData    => PPCDMDCRDBUSOUT8_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(8)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(8),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(8),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(9),
	GlitchData    => PPCDMDCRDBUSOUT9_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(9)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(9),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(9),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(10),
	GlitchData    => PPCDMDCRDBUSOUT10_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(10)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(10),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(10),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(11),
	GlitchData    => PPCDMDCRDBUSOUT11_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(11)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(11),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(11),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(12),
	GlitchData    => PPCDMDCRDBUSOUT12_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(12)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(12),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(12),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(13),
	GlitchData    => PPCDMDCRDBUSOUT13_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(13)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(13),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(13),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(14),
	GlitchData    => PPCDMDCRDBUSOUT14_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(14)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(14),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(14),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(15),
	GlitchData    => PPCDMDCRDBUSOUT15_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(15)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(15),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(15),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(16),
	GlitchData    => PPCDMDCRDBUSOUT16_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(16)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(16),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(16),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(17),
	GlitchData    => PPCDMDCRDBUSOUT17_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(17)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(17),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(17),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(18),
	GlitchData    => PPCDMDCRDBUSOUT18_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(18)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(18),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(18),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(19),
	GlitchData    => PPCDMDCRDBUSOUT19_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(19)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(19),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(19),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(20),
	GlitchData    => PPCDMDCRDBUSOUT20_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(20)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(20),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(20),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(21),
	GlitchData    => PPCDMDCRDBUSOUT21_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(21)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(21),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(21),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(22),
	GlitchData    => PPCDMDCRDBUSOUT22_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(22)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(22),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(22),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(23),
	GlitchData    => PPCDMDCRDBUSOUT23_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(23)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(23),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(23),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(24),
	GlitchData    => PPCDMDCRDBUSOUT24_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(24)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(24),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(24),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(25),
	GlitchData    => PPCDMDCRDBUSOUT25_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(25)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(25),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(25),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(26),
	GlitchData    => PPCDMDCRDBUSOUT26_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(26)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(26),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(26),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(27),
	GlitchData    => PPCDMDCRDBUSOUT27_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(27)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(27),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(27),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(28),
	GlitchData    => PPCDMDCRDBUSOUT28_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(28)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(28),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(28),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(29),
	GlitchData    => PPCDMDCRDBUSOUT29_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(29)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(29),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(29),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(30),
	GlitchData    => PPCDMDCRDBUSOUT30_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(30)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(30),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(30),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRDBUSOUT(31),
	GlitchData    => PPCDMDCRDBUSOUT31_GlitchData,
	OutSignalName => "PPCDMDCRDBUSOUT(31)",
	OutTemp       => PPCDMDCRDBUSOUT_OUT(31),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(31),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRDBUSOUT(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRREAD,
	GlitchData    => PPCDMDCRREAD_GlitchData,
	OutSignalName => "PPCDMDCRREAD",
	OutTemp       => PPCDMDCRREAD_OUT,
	Paths         => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRREAD,TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRREAD, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRUABUS(20),
	GlitchData    => PPCDMDCRUABUS20_GlitchData,
	OutSignalName => "PPCDMDCRUABUS(20)",
	OutTemp       => PPCDMDCRUABUS_OUT(20),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRUABUS(20),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRUABUS(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRUABUS(21),
	GlitchData    => PPCDMDCRUABUS21_GlitchData,
	OutSignalName => "PPCDMDCRUABUS(21)",
	OutTemp       => PPCDMDCRUABUS_OUT(21),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRUABUS(21),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRUABUS(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDMDCRWRITE,
	GlitchData    => PPCDMDCRWRITE_GlitchData,
	OutSignalName => "PPCDMDCRWRITE",
	OutTemp       => PPCDMDCRWRITE_OUT,
	Paths         => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDMDCRWRITE,TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDMDCRWRITE, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABORT,
	GlitchData    => PPCMPLBABORT_GlitchData,
	OutSignalName => "PPCMPLBABORT",
	OutTemp       => PPCMPLBABORT_OUT,
	Paths         => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABORT,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABORT, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(0),
	GlitchData    => PPCMPLBABUS0_GlitchData,
	OutSignalName => "PPCMPLBABUS(0)",
	OutTemp       => PPCMPLBABUS_OUT(0),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(1),
	GlitchData    => PPCMPLBABUS1_GlitchData,
	OutSignalName => "PPCMPLBABUS(1)",
	OutTemp       => PPCMPLBABUS_OUT(1),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(2),
	GlitchData    => PPCMPLBABUS2_GlitchData,
	OutSignalName => "PPCMPLBABUS(2)",
	OutTemp       => PPCMPLBABUS_OUT(2),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(3),
	GlitchData    => PPCMPLBABUS3_GlitchData,
	OutSignalName => "PPCMPLBABUS(3)",
	OutTemp       => PPCMPLBABUS_OUT(3),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(4),
	GlitchData    => PPCMPLBABUS4_GlitchData,
	OutSignalName => "PPCMPLBABUS(4)",
	OutTemp       => PPCMPLBABUS_OUT(4),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(4),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(5),
	GlitchData    => PPCMPLBABUS5_GlitchData,
	OutSignalName => "PPCMPLBABUS(5)",
	OutTemp       => PPCMPLBABUS_OUT(5),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(5),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(6),
	GlitchData    => PPCMPLBABUS6_GlitchData,
	OutSignalName => "PPCMPLBABUS(6)",
	OutTemp       => PPCMPLBABUS_OUT(6),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(6),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(7),
	GlitchData    => PPCMPLBABUS7_GlitchData,
	OutSignalName => "PPCMPLBABUS(7)",
	OutTemp       => PPCMPLBABUS_OUT(7),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(7),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(8),
	GlitchData    => PPCMPLBABUS8_GlitchData,
	OutSignalName => "PPCMPLBABUS(8)",
	OutTemp       => PPCMPLBABUS_OUT(8),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(8),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(9),
	GlitchData    => PPCMPLBABUS9_GlitchData,
	OutSignalName => "PPCMPLBABUS(9)",
	OutTemp       => PPCMPLBABUS_OUT(9),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(9),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(10),
	GlitchData    => PPCMPLBABUS10_GlitchData,
	OutSignalName => "PPCMPLBABUS(10)",
	OutTemp       => PPCMPLBABUS_OUT(10),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(10),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(11),
	GlitchData    => PPCMPLBABUS11_GlitchData,
	OutSignalName => "PPCMPLBABUS(11)",
	OutTemp       => PPCMPLBABUS_OUT(11),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(11),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(12),
	GlitchData    => PPCMPLBABUS12_GlitchData,
	OutSignalName => "PPCMPLBABUS(12)",
	OutTemp       => PPCMPLBABUS_OUT(12),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(12),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(13),
	GlitchData    => PPCMPLBABUS13_GlitchData,
	OutSignalName => "PPCMPLBABUS(13)",
	OutTemp       => PPCMPLBABUS_OUT(13),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(13),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(14),
	GlitchData    => PPCMPLBABUS14_GlitchData,
	OutSignalName => "PPCMPLBABUS(14)",
	OutTemp       => PPCMPLBABUS_OUT(14),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(14),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(15),
	GlitchData    => PPCMPLBABUS15_GlitchData,
	OutSignalName => "PPCMPLBABUS(15)",
	OutTemp       => PPCMPLBABUS_OUT(15),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(15),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(16),
	GlitchData    => PPCMPLBABUS16_GlitchData,
	OutSignalName => "PPCMPLBABUS(16)",
	OutTemp       => PPCMPLBABUS_OUT(16),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(16),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(17),
	GlitchData    => PPCMPLBABUS17_GlitchData,
	OutSignalName => "PPCMPLBABUS(17)",
	OutTemp       => PPCMPLBABUS_OUT(17),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(17),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(18),
	GlitchData    => PPCMPLBABUS18_GlitchData,
	OutSignalName => "PPCMPLBABUS(18)",
	OutTemp       => PPCMPLBABUS_OUT(18),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(18),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(19),
	GlitchData    => PPCMPLBABUS19_GlitchData,
	OutSignalName => "PPCMPLBABUS(19)",
	OutTemp       => PPCMPLBABUS_OUT(19),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(19),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(20),
	GlitchData    => PPCMPLBABUS20_GlitchData,
	OutSignalName => "PPCMPLBABUS(20)",
	OutTemp       => PPCMPLBABUS_OUT(20),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(20),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(21),
	GlitchData    => PPCMPLBABUS21_GlitchData,
	OutSignalName => "PPCMPLBABUS(21)",
	OutTemp       => PPCMPLBABUS_OUT(21),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(21),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(22),
	GlitchData    => PPCMPLBABUS22_GlitchData,
	OutSignalName => "PPCMPLBABUS(22)",
	OutTemp       => PPCMPLBABUS_OUT(22),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(22),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(23),
	GlitchData    => PPCMPLBABUS23_GlitchData,
	OutSignalName => "PPCMPLBABUS(23)",
	OutTemp       => PPCMPLBABUS_OUT(23),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(23),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(24),
	GlitchData    => PPCMPLBABUS24_GlitchData,
	OutSignalName => "PPCMPLBABUS(24)",
	OutTemp       => PPCMPLBABUS_OUT(24),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(24),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(25),
	GlitchData    => PPCMPLBABUS25_GlitchData,
	OutSignalName => "PPCMPLBABUS(25)",
	OutTemp       => PPCMPLBABUS_OUT(25),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(25),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(26),
	GlitchData    => PPCMPLBABUS26_GlitchData,
	OutSignalName => "PPCMPLBABUS(26)",
	OutTemp       => PPCMPLBABUS_OUT(26),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(26),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(27),
	GlitchData    => PPCMPLBABUS27_GlitchData,
	OutSignalName => "PPCMPLBABUS(27)",
	OutTemp       => PPCMPLBABUS_OUT(27),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(27),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(28),
	GlitchData    => PPCMPLBABUS28_GlitchData,
	OutSignalName => "PPCMPLBABUS(28)",
	OutTemp       => PPCMPLBABUS_OUT(28),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(28),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(29),
	GlitchData    => PPCMPLBABUS29_GlitchData,
	OutSignalName => "PPCMPLBABUS(29)",
	OutTemp       => PPCMPLBABUS_OUT(29),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(29),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(30),
	GlitchData    => PPCMPLBABUS30_GlitchData,
	OutSignalName => "PPCMPLBABUS(30)",
	OutTemp       => PPCMPLBABUS_OUT(30),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(30),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBABUS(31),
	GlitchData    => PPCMPLBABUS31_GlitchData,
	OutSignalName => "PPCMPLBABUS(31)",
	OutTemp       => PPCMPLBABUS_OUT(31),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBABUS(31),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBABUS(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(0),
	GlitchData    => PPCMPLBBE0_GlitchData,
	OutSignalName => "PPCMPLBBE(0)",
	OutTemp       => PPCMPLBBE_OUT(0),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(1),
	GlitchData    => PPCMPLBBE1_GlitchData,
	OutSignalName => "PPCMPLBBE(1)",
	OutTemp       => PPCMPLBBE_OUT(1),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(2),
	GlitchData    => PPCMPLBBE2_GlitchData,
	OutSignalName => "PPCMPLBBE(2)",
	OutTemp       => PPCMPLBBE_OUT(2),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(3),
	GlitchData    => PPCMPLBBE3_GlitchData,
	OutSignalName => "PPCMPLBBE(3)",
	OutTemp       => PPCMPLBBE_OUT(3),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(4),
	GlitchData    => PPCMPLBBE4_GlitchData,
	OutSignalName => "PPCMPLBBE(4)",
	OutTemp       => PPCMPLBBE_OUT(4),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(4),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(5),
	GlitchData    => PPCMPLBBE5_GlitchData,
	OutSignalName => "PPCMPLBBE(5)",
	OutTemp       => PPCMPLBBE_OUT(5),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(5),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(6),
	GlitchData    => PPCMPLBBE6_GlitchData,
	OutSignalName => "PPCMPLBBE(6)",
	OutTemp       => PPCMPLBBE_OUT(6),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(6),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(7),
	GlitchData    => PPCMPLBBE7_GlitchData,
	OutSignalName => "PPCMPLBBE(7)",
	OutTemp       => PPCMPLBBE_OUT(7),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(7),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(8),
	GlitchData    => PPCMPLBBE8_GlitchData,
	OutSignalName => "PPCMPLBBE(8)",
	OutTemp       => PPCMPLBBE_OUT(8),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(8),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(9),
	GlitchData    => PPCMPLBBE9_GlitchData,
	OutSignalName => "PPCMPLBBE(9)",
	OutTemp       => PPCMPLBBE_OUT(9),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(9),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(10),
	GlitchData    => PPCMPLBBE10_GlitchData,
	OutSignalName => "PPCMPLBBE(10)",
	OutTemp       => PPCMPLBBE_OUT(10),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(10),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(11),
	GlitchData    => PPCMPLBBE11_GlitchData,
	OutSignalName => "PPCMPLBBE(11)",
	OutTemp       => PPCMPLBBE_OUT(11),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(11),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(12),
	GlitchData    => PPCMPLBBE12_GlitchData,
	OutSignalName => "PPCMPLBBE(12)",
	OutTemp       => PPCMPLBBE_OUT(12),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(12),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(13),
	GlitchData    => PPCMPLBBE13_GlitchData,
	OutSignalName => "PPCMPLBBE(13)",
	OutTemp       => PPCMPLBBE_OUT(13),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(13),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(14),
	GlitchData    => PPCMPLBBE14_GlitchData,
	OutSignalName => "PPCMPLBBE(14)",
	OutTemp       => PPCMPLBBE_OUT(14),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(14),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBE(15),
	GlitchData    => PPCMPLBBE15_GlitchData,
	OutSignalName => "PPCMPLBBE(15)",
	OutTemp       => PPCMPLBBE_OUT(15),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBE(15),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBE(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBBUSLOCK,
	GlitchData    => PPCMPLBBUSLOCK_GlitchData,
	OutSignalName => "PPCMPLBBUSLOCK",
	OutTemp       => PPCMPLBBUSLOCK_OUT,
	Paths         => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBBUSLOCK,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBBUSLOCK, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBLOCKERR,
	GlitchData    => PPCMPLBLOCKERR_GlitchData,
	OutSignalName => "PPCMPLBLOCKERR",
	OutTemp       => PPCMPLBLOCKERR_OUT,
	Paths         => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBLOCKERR,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBLOCKERR, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBPRIORITY(0),
	GlitchData    => PPCMPLBPRIORITY0_GlitchData,
	OutSignalName => "PPCMPLBPRIORITY(0)",
	OutTemp       => PPCMPLBPRIORITY_OUT(0),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBPRIORITY(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBPRIORITY(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBPRIORITY(1),
	GlitchData    => PPCMPLBPRIORITY1_GlitchData,
	OutSignalName => "PPCMPLBPRIORITY(1)",
	OutTemp       => PPCMPLBPRIORITY_OUT(1),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBPRIORITY(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBPRIORITY(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBRDBURST,
	GlitchData    => PPCMPLBRDBURST_GlitchData,
	OutSignalName => "PPCMPLBRDBURST",
	OutTemp       => PPCMPLBRDBURST_OUT,
	Paths         => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBRDBURST,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBRDBURST, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBREQUEST,
	GlitchData    => PPCMPLBREQUEST_GlitchData,
	OutSignalName => "PPCMPLBREQUEST",
	OutTemp       => PPCMPLBREQUEST_OUT,
	Paths         => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBREQUEST,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBREQUEST, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBRNW,
	GlitchData    => PPCMPLBRNW_GlitchData,
	OutSignalName => "PPCMPLBRNW",
	OutTemp       => PPCMPLBRNW_OUT,
	Paths         => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBRNW,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBRNW, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBSIZE(0),
	GlitchData    => PPCMPLBSIZE0_GlitchData,
	OutSignalName => "PPCMPLBSIZE(0)",
	OutTemp       => PPCMPLBSIZE_OUT(0),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBSIZE(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBSIZE(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBSIZE(1),
	GlitchData    => PPCMPLBSIZE1_GlitchData,
	OutSignalName => "PPCMPLBSIZE(1)",
	OutTemp       => PPCMPLBSIZE_OUT(1),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBSIZE(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBSIZE(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBSIZE(2),
	GlitchData    => PPCMPLBSIZE2_GlitchData,
	OutSignalName => "PPCMPLBSIZE(2)",
	OutTemp       => PPCMPLBSIZE_OUT(2),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBSIZE(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBSIZE(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBSIZE(3),
	GlitchData    => PPCMPLBSIZE3_GlitchData,
	OutSignalName => "PPCMPLBSIZE(3)",
	OutTemp       => PPCMPLBSIZE_OUT(3),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBSIZE(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBSIZE(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(0),
	GlitchData    => PPCMPLBTATTRIBUTE0_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(0)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(0),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(1),
	GlitchData    => PPCMPLBTATTRIBUTE1_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(1)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(1),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(2),
	GlitchData    => PPCMPLBTATTRIBUTE2_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(2)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(2),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(3),
	GlitchData    => PPCMPLBTATTRIBUTE3_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(3)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(3),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(4),
	GlitchData    => PPCMPLBTATTRIBUTE4_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(4)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(4),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(4),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(5),
	GlitchData    => PPCMPLBTATTRIBUTE5_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(5)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(5),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(5),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(6),
	GlitchData    => PPCMPLBTATTRIBUTE6_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(6)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(6),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(6),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(7),
	GlitchData    => PPCMPLBTATTRIBUTE7_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(7)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(7),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(7),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(8),
	GlitchData    => PPCMPLBTATTRIBUTE8_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(8)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(8),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(8),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(9),
	GlitchData    => PPCMPLBTATTRIBUTE9_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(9)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(9),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(9),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(10),
	GlitchData    => PPCMPLBTATTRIBUTE10_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(10)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(10),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(10),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(11),
	GlitchData    => PPCMPLBTATTRIBUTE11_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(11)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(11),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(11),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(12),
	GlitchData    => PPCMPLBTATTRIBUTE12_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(12)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(12),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(12),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(13),
	GlitchData    => PPCMPLBTATTRIBUTE13_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(13)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(13),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(13),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(14),
	GlitchData    => PPCMPLBTATTRIBUTE14_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(14)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(14),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(14),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTATTRIBUTE(15),
	GlitchData    => PPCMPLBTATTRIBUTE15_GlitchData,
	OutSignalName => "PPCMPLBTATTRIBUTE(15)",
	OutTemp       => PPCMPLBTATTRIBUTE_OUT(15),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(15),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTATTRIBUTE(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTYPE(0),
	GlitchData    => PPCMPLBTYPE0_GlitchData,
	OutSignalName => "PPCMPLBTYPE(0)",
	OutTemp       => PPCMPLBTYPE_OUT(0),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTYPE(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTYPE(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTYPE(1),
	GlitchData    => PPCMPLBTYPE1_GlitchData,
	OutSignalName => "PPCMPLBTYPE(1)",
	OutTemp       => PPCMPLBTYPE_OUT(1),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTYPE(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTYPE(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBTYPE(2),
	GlitchData    => PPCMPLBTYPE2_GlitchData,
	OutSignalName => "PPCMPLBTYPE(2)",
	OutTemp       => PPCMPLBTYPE_OUT(2),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBTYPE(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBTYPE(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBUABUS(28),
	GlitchData    => PPCMPLBUABUS28_GlitchData,
	OutSignalName => "PPCMPLBUABUS(28)",
	OutTemp       => PPCMPLBUABUS_OUT(28),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBUABUS(28),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBUABUS(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBUABUS(29),
	GlitchData    => PPCMPLBUABUS29_GlitchData,
	OutSignalName => "PPCMPLBUABUS(29)",
	OutTemp       => PPCMPLBUABUS_OUT(29),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBUABUS(29),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBUABUS(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBUABUS(30),
	GlitchData    => PPCMPLBUABUS30_GlitchData,
	OutSignalName => "PPCMPLBUABUS(30)",
	OutTemp       => PPCMPLBUABUS_OUT(30),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBUABUS(30),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBUABUS(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBUABUS(31),
	GlitchData    => PPCMPLBUABUS31_GlitchData,
	OutSignalName => "PPCMPLBUABUS(31)",
	OutTemp       => PPCMPLBUABUS_OUT(31),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBUABUS(31),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBUABUS(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRBURST,
	GlitchData    => PPCMPLBWRBURST_GlitchData,
	OutSignalName => "PPCMPLBWRBURST",
	OutTemp       => PPCMPLBWRBURST_OUT,
	Paths         => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRBURST,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRBURST, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(0),
	GlitchData    => PPCMPLBWRDBUS0_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(0)",
	OutTemp       => PPCMPLBWRDBUS_OUT(0),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(1),
	GlitchData    => PPCMPLBWRDBUS1_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(1)",
	OutTemp       => PPCMPLBWRDBUS_OUT(1),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(2),
	GlitchData    => PPCMPLBWRDBUS2_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(2)",
	OutTemp       => PPCMPLBWRDBUS_OUT(2),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(3),
	GlitchData    => PPCMPLBWRDBUS3_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(3)",
	OutTemp       => PPCMPLBWRDBUS_OUT(3),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(4),
	GlitchData    => PPCMPLBWRDBUS4_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(4)",
	OutTemp       => PPCMPLBWRDBUS_OUT(4),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(4),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(5),
	GlitchData    => PPCMPLBWRDBUS5_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(5)",
	OutTemp       => PPCMPLBWRDBUS_OUT(5),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(5),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(6),
	GlitchData    => PPCMPLBWRDBUS6_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(6)",
	OutTemp       => PPCMPLBWRDBUS_OUT(6),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(6),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(7),
	GlitchData    => PPCMPLBWRDBUS7_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(7)",
	OutTemp       => PPCMPLBWRDBUS_OUT(7),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(7),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(8),
	GlitchData    => PPCMPLBWRDBUS8_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(8)",
	OutTemp       => PPCMPLBWRDBUS_OUT(8),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(8),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(9),
	GlitchData    => PPCMPLBWRDBUS9_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(9)",
	OutTemp       => PPCMPLBWRDBUS_OUT(9),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(9),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(10),
	GlitchData    => PPCMPLBWRDBUS10_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(10)",
	OutTemp       => PPCMPLBWRDBUS_OUT(10),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(10),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(11),
	GlitchData    => PPCMPLBWRDBUS11_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(11)",
	OutTemp       => PPCMPLBWRDBUS_OUT(11),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(11),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(12),
	GlitchData    => PPCMPLBWRDBUS12_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(12)",
	OutTemp       => PPCMPLBWRDBUS_OUT(12),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(12),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(13),
	GlitchData    => PPCMPLBWRDBUS13_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(13)",
	OutTemp       => PPCMPLBWRDBUS_OUT(13),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(13),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(14),
	GlitchData    => PPCMPLBWRDBUS14_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(14)",
	OutTemp       => PPCMPLBWRDBUS_OUT(14),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(14),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(15),
	GlitchData    => PPCMPLBWRDBUS15_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(15)",
	OutTemp       => PPCMPLBWRDBUS_OUT(15),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(15),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(16),
	GlitchData    => PPCMPLBWRDBUS16_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(16)",
	OutTemp       => PPCMPLBWRDBUS_OUT(16),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(16),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(17),
	GlitchData    => PPCMPLBWRDBUS17_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(17)",
	OutTemp       => PPCMPLBWRDBUS_OUT(17),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(17),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(18),
	GlitchData    => PPCMPLBWRDBUS18_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(18)",
	OutTemp       => PPCMPLBWRDBUS_OUT(18),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(18),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(19),
	GlitchData    => PPCMPLBWRDBUS19_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(19)",
	OutTemp       => PPCMPLBWRDBUS_OUT(19),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(19),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(20),
	GlitchData    => PPCMPLBWRDBUS20_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(20)",
	OutTemp       => PPCMPLBWRDBUS_OUT(20),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(20),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(21),
	GlitchData    => PPCMPLBWRDBUS21_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(21)",
	OutTemp       => PPCMPLBWRDBUS_OUT(21),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(21),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(22),
	GlitchData    => PPCMPLBWRDBUS22_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(22)",
	OutTemp       => PPCMPLBWRDBUS_OUT(22),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(22),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(23),
	GlitchData    => PPCMPLBWRDBUS23_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(23)",
	OutTemp       => PPCMPLBWRDBUS_OUT(23),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(23),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(24),
	GlitchData    => PPCMPLBWRDBUS24_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(24)",
	OutTemp       => PPCMPLBWRDBUS_OUT(24),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(24),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(25),
	GlitchData    => PPCMPLBWRDBUS25_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(25)",
	OutTemp       => PPCMPLBWRDBUS_OUT(25),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(25),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(26),
	GlitchData    => PPCMPLBWRDBUS26_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(26)",
	OutTemp       => PPCMPLBWRDBUS_OUT(26),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(26),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(27),
	GlitchData    => PPCMPLBWRDBUS27_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(27)",
	OutTemp       => PPCMPLBWRDBUS_OUT(27),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(27),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(28),
	GlitchData    => PPCMPLBWRDBUS28_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(28)",
	OutTemp       => PPCMPLBWRDBUS_OUT(28),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(28),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(29),
	GlitchData    => PPCMPLBWRDBUS29_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(29)",
	OutTemp       => PPCMPLBWRDBUS_OUT(29),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(29),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(30),
	GlitchData    => PPCMPLBWRDBUS30_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(30)",
	OutTemp       => PPCMPLBWRDBUS_OUT(30),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(30),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(31),
	GlitchData    => PPCMPLBWRDBUS31_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(31)",
	OutTemp       => PPCMPLBWRDBUS_OUT(31),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(31),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(32),
	GlitchData    => PPCMPLBWRDBUS32_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(32)",
	OutTemp       => PPCMPLBWRDBUS_OUT(32),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(32),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(32), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(33),
	GlitchData    => PPCMPLBWRDBUS33_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(33)",
	OutTemp       => PPCMPLBWRDBUS_OUT(33),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(33),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(33), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(34),
	GlitchData    => PPCMPLBWRDBUS34_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(34)",
	OutTemp       => PPCMPLBWRDBUS_OUT(34),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(34),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(34), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(35),
	GlitchData    => PPCMPLBWRDBUS35_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(35)",
	OutTemp       => PPCMPLBWRDBUS_OUT(35),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(35),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(35), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(36),
	GlitchData    => PPCMPLBWRDBUS36_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(36)",
	OutTemp       => PPCMPLBWRDBUS_OUT(36),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(36),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(36), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(37),
	GlitchData    => PPCMPLBWRDBUS37_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(37)",
	OutTemp       => PPCMPLBWRDBUS_OUT(37),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(37),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(37), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(38),
	GlitchData    => PPCMPLBWRDBUS38_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(38)",
	OutTemp       => PPCMPLBWRDBUS_OUT(38),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(38),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(38), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(39),
	GlitchData    => PPCMPLBWRDBUS39_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(39)",
	OutTemp       => PPCMPLBWRDBUS_OUT(39),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(39),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(39), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(40),
	GlitchData    => PPCMPLBWRDBUS40_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(40)",
	OutTemp       => PPCMPLBWRDBUS_OUT(40),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(40),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(40), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(41),
	GlitchData    => PPCMPLBWRDBUS41_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(41)",
	OutTemp       => PPCMPLBWRDBUS_OUT(41),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(41),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(41), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(42),
	GlitchData    => PPCMPLBWRDBUS42_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(42)",
	OutTemp       => PPCMPLBWRDBUS_OUT(42),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(42),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(42), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(43),
	GlitchData    => PPCMPLBWRDBUS43_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(43)",
	OutTemp       => PPCMPLBWRDBUS_OUT(43),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(43),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(43), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(44),
	GlitchData    => PPCMPLBWRDBUS44_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(44)",
	OutTemp       => PPCMPLBWRDBUS_OUT(44),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(44),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(44), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(45),
	GlitchData    => PPCMPLBWRDBUS45_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(45)",
	OutTemp       => PPCMPLBWRDBUS_OUT(45),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(45),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(45), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(46),
	GlitchData    => PPCMPLBWRDBUS46_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(46)",
	OutTemp       => PPCMPLBWRDBUS_OUT(46),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(46),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(46), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(47),
	GlitchData    => PPCMPLBWRDBUS47_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(47)",
	OutTemp       => PPCMPLBWRDBUS_OUT(47),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(47),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(47), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(48),
	GlitchData    => PPCMPLBWRDBUS48_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(48)",
	OutTemp       => PPCMPLBWRDBUS_OUT(48),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(48),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(48), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(49),
	GlitchData    => PPCMPLBWRDBUS49_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(49)",
	OutTemp       => PPCMPLBWRDBUS_OUT(49),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(49),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(49), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(50),
	GlitchData    => PPCMPLBWRDBUS50_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(50)",
	OutTemp       => PPCMPLBWRDBUS_OUT(50),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(50),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(50), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(51),
	GlitchData    => PPCMPLBWRDBUS51_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(51)",
	OutTemp       => PPCMPLBWRDBUS_OUT(51),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(51),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(51), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(52),
	GlitchData    => PPCMPLBWRDBUS52_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(52)",
	OutTemp       => PPCMPLBWRDBUS_OUT(52),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(52),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(52), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(53),
	GlitchData    => PPCMPLBWRDBUS53_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(53)",
	OutTemp       => PPCMPLBWRDBUS_OUT(53),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(53),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(53), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(54),
	GlitchData    => PPCMPLBWRDBUS54_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(54)",
	OutTemp       => PPCMPLBWRDBUS_OUT(54),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(54),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(54), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(55),
	GlitchData    => PPCMPLBWRDBUS55_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(55)",
	OutTemp       => PPCMPLBWRDBUS_OUT(55),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(55),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(55), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(56),
	GlitchData    => PPCMPLBWRDBUS56_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(56)",
	OutTemp       => PPCMPLBWRDBUS_OUT(56),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(56),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(56), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(57),
	GlitchData    => PPCMPLBWRDBUS57_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(57)",
	OutTemp       => PPCMPLBWRDBUS_OUT(57),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(57),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(57), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(58),
	GlitchData    => PPCMPLBWRDBUS58_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(58)",
	OutTemp       => PPCMPLBWRDBUS_OUT(58),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(58),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(58), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(59),
	GlitchData    => PPCMPLBWRDBUS59_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(59)",
	OutTemp       => PPCMPLBWRDBUS_OUT(59),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(59),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(59), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(60),
	GlitchData    => PPCMPLBWRDBUS60_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(60)",
	OutTemp       => PPCMPLBWRDBUS_OUT(60),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(60),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(60), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(61),
	GlitchData    => PPCMPLBWRDBUS61_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(61)",
	OutTemp       => PPCMPLBWRDBUS_OUT(61),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(61),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(61), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(62),
	GlitchData    => PPCMPLBWRDBUS62_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(62)",
	OutTemp       => PPCMPLBWRDBUS_OUT(62),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(62),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(62), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(63),
	GlitchData    => PPCMPLBWRDBUS63_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(63)",
	OutTemp       => PPCMPLBWRDBUS_OUT(63),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(63),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(63), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(64),
	GlitchData    => PPCMPLBWRDBUS64_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(64)",
	OutTemp       => PPCMPLBWRDBUS_OUT(64),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(64),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(64), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(65),
	GlitchData    => PPCMPLBWRDBUS65_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(65)",
	OutTemp       => PPCMPLBWRDBUS_OUT(65),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(65),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(65), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(66),
	GlitchData    => PPCMPLBWRDBUS66_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(66)",
	OutTemp       => PPCMPLBWRDBUS_OUT(66),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(66),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(66), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(67),
	GlitchData    => PPCMPLBWRDBUS67_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(67)",
	OutTemp       => PPCMPLBWRDBUS_OUT(67),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(67),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(67), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(68),
	GlitchData    => PPCMPLBWRDBUS68_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(68)",
	OutTemp       => PPCMPLBWRDBUS_OUT(68),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(68),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(68), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(69),
	GlitchData    => PPCMPLBWRDBUS69_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(69)",
	OutTemp       => PPCMPLBWRDBUS_OUT(69),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(69),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(69), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(70),
	GlitchData    => PPCMPLBWRDBUS70_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(70)",
	OutTemp       => PPCMPLBWRDBUS_OUT(70),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(70),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(70), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(71),
	GlitchData    => PPCMPLBWRDBUS71_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(71)",
	OutTemp       => PPCMPLBWRDBUS_OUT(71),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(71),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(71), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(72),
	GlitchData    => PPCMPLBWRDBUS72_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(72)",
	OutTemp       => PPCMPLBWRDBUS_OUT(72),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(72),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(72), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(73),
	GlitchData    => PPCMPLBWRDBUS73_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(73)",
	OutTemp       => PPCMPLBWRDBUS_OUT(73),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(73),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(73), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(74),
	GlitchData    => PPCMPLBWRDBUS74_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(74)",
	OutTemp       => PPCMPLBWRDBUS_OUT(74),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(74),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(74), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(75),
	GlitchData    => PPCMPLBWRDBUS75_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(75)",
	OutTemp       => PPCMPLBWRDBUS_OUT(75),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(75),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(75), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(76),
	GlitchData    => PPCMPLBWRDBUS76_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(76)",
	OutTemp       => PPCMPLBWRDBUS_OUT(76),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(76),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(76), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(77),
	GlitchData    => PPCMPLBWRDBUS77_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(77)",
	OutTemp       => PPCMPLBWRDBUS_OUT(77),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(77),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(77), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(78),
	GlitchData    => PPCMPLBWRDBUS78_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(78)",
	OutTemp       => PPCMPLBWRDBUS_OUT(78),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(78),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(78), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(79),
	GlitchData    => PPCMPLBWRDBUS79_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(79)",
	OutTemp       => PPCMPLBWRDBUS_OUT(79),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(79),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(79), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(80),
	GlitchData    => PPCMPLBWRDBUS80_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(80)",
	OutTemp       => PPCMPLBWRDBUS_OUT(80),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(80),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(80), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(81),
	GlitchData    => PPCMPLBWRDBUS81_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(81)",
	OutTemp       => PPCMPLBWRDBUS_OUT(81),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(81),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(81), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(82),
	GlitchData    => PPCMPLBWRDBUS82_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(82)",
	OutTemp       => PPCMPLBWRDBUS_OUT(82),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(82),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(82), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(83),
	GlitchData    => PPCMPLBWRDBUS83_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(83)",
	OutTemp       => PPCMPLBWRDBUS_OUT(83),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(83),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(83), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(84),
	GlitchData    => PPCMPLBWRDBUS84_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(84)",
	OutTemp       => PPCMPLBWRDBUS_OUT(84),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(84),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(84), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(85),
	GlitchData    => PPCMPLBWRDBUS85_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(85)",
	OutTemp       => PPCMPLBWRDBUS_OUT(85),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(85),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(85), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(86),
	GlitchData    => PPCMPLBWRDBUS86_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(86)",
	OutTemp       => PPCMPLBWRDBUS_OUT(86),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(86),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(86), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(87),
	GlitchData    => PPCMPLBWRDBUS87_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(87)",
	OutTemp       => PPCMPLBWRDBUS_OUT(87),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(87),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(87), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(88),
	GlitchData    => PPCMPLBWRDBUS88_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(88)",
	OutTemp       => PPCMPLBWRDBUS_OUT(88),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(88),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(88), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(89),
	GlitchData    => PPCMPLBWRDBUS89_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(89)",
	OutTemp       => PPCMPLBWRDBUS_OUT(89),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(89),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(89), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(90),
	GlitchData    => PPCMPLBWRDBUS90_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(90)",
	OutTemp       => PPCMPLBWRDBUS_OUT(90),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(90),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(90), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(91),
	GlitchData    => PPCMPLBWRDBUS91_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(91)",
	OutTemp       => PPCMPLBWRDBUS_OUT(91),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(91),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(91), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(92),
	GlitchData    => PPCMPLBWRDBUS92_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(92)",
	OutTemp       => PPCMPLBWRDBUS_OUT(92),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(92),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(92), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(93),
	GlitchData    => PPCMPLBWRDBUS93_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(93)",
	OutTemp       => PPCMPLBWRDBUS_OUT(93),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(93),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(93), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(94),
	GlitchData    => PPCMPLBWRDBUS94_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(94)",
	OutTemp       => PPCMPLBWRDBUS_OUT(94),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(94),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(94), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(95),
	GlitchData    => PPCMPLBWRDBUS95_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(95)",
	OutTemp       => PPCMPLBWRDBUS_OUT(95),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(95),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(95), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(96),
	GlitchData    => PPCMPLBWRDBUS96_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(96)",
	OutTemp       => PPCMPLBWRDBUS_OUT(96),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(96),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(96), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(97),
	GlitchData    => PPCMPLBWRDBUS97_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(97)",
	OutTemp       => PPCMPLBWRDBUS_OUT(97),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(97),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(97), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(98),
	GlitchData    => PPCMPLBWRDBUS98_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(98)",
	OutTemp       => PPCMPLBWRDBUS_OUT(98),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(98),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(98), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(99),
	GlitchData    => PPCMPLBWRDBUS99_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(99)",
	OutTemp       => PPCMPLBWRDBUS_OUT(99),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(99),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(99), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(100),
	GlitchData    => PPCMPLBWRDBUS100_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(100)",
	OutTemp       => PPCMPLBWRDBUS_OUT(100),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(100),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(100), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(101),
	GlitchData    => PPCMPLBWRDBUS101_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(101)",
	OutTemp       => PPCMPLBWRDBUS_OUT(101),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(101),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(101), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(102),
	GlitchData    => PPCMPLBWRDBUS102_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(102)",
	OutTemp       => PPCMPLBWRDBUS_OUT(102),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(102),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(102), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(103),
	GlitchData    => PPCMPLBWRDBUS103_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(103)",
	OutTemp       => PPCMPLBWRDBUS_OUT(103),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(103),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(103), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(104),
	GlitchData    => PPCMPLBWRDBUS104_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(104)",
	OutTemp       => PPCMPLBWRDBUS_OUT(104),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(104),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(104), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(105),
	GlitchData    => PPCMPLBWRDBUS105_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(105)",
	OutTemp       => PPCMPLBWRDBUS_OUT(105),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(105),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(105), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(106),
	GlitchData    => PPCMPLBWRDBUS106_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(106)",
	OutTemp       => PPCMPLBWRDBUS_OUT(106),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(106),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(106), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(107),
	GlitchData    => PPCMPLBWRDBUS107_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(107)",
	OutTemp       => PPCMPLBWRDBUS_OUT(107),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(107),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(107), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(108),
	GlitchData    => PPCMPLBWRDBUS108_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(108)",
	OutTemp       => PPCMPLBWRDBUS_OUT(108),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(108),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(108), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(109),
	GlitchData    => PPCMPLBWRDBUS109_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(109)",
	OutTemp       => PPCMPLBWRDBUS_OUT(109),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(109),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(109), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(110),
	GlitchData    => PPCMPLBWRDBUS110_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(110)",
	OutTemp       => PPCMPLBWRDBUS_OUT(110),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(110),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(110), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(111),
	GlitchData    => PPCMPLBWRDBUS111_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(111)",
	OutTemp       => PPCMPLBWRDBUS_OUT(111),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(111),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(111), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(112),
	GlitchData    => PPCMPLBWRDBUS112_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(112)",
	OutTemp       => PPCMPLBWRDBUS_OUT(112),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(112),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(112), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(113),
	GlitchData    => PPCMPLBWRDBUS113_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(113)",
	OutTemp       => PPCMPLBWRDBUS_OUT(113),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(113),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(113), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(114),
	GlitchData    => PPCMPLBWRDBUS114_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(114)",
	OutTemp       => PPCMPLBWRDBUS_OUT(114),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(114),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(114), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(115),
	GlitchData    => PPCMPLBWRDBUS115_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(115)",
	OutTemp       => PPCMPLBWRDBUS_OUT(115),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(115),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(115), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(116),
	GlitchData    => PPCMPLBWRDBUS116_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(116)",
	OutTemp       => PPCMPLBWRDBUS_OUT(116),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(116),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(116), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(117),
	GlitchData    => PPCMPLBWRDBUS117_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(117)",
	OutTemp       => PPCMPLBWRDBUS_OUT(117),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(117),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(117), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(118),
	GlitchData    => PPCMPLBWRDBUS118_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(118)",
	OutTemp       => PPCMPLBWRDBUS_OUT(118),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(118),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(118), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(119),
	GlitchData    => PPCMPLBWRDBUS119_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(119)",
	OutTemp       => PPCMPLBWRDBUS_OUT(119),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(119),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(119), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(120),
	GlitchData    => PPCMPLBWRDBUS120_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(120)",
	OutTemp       => PPCMPLBWRDBUS_OUT(120),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(120),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(120), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(121),
	GlitchData    => PPCMPLBWRDBUS121_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(121)",
	OutTemp       => PPCMPLBWRDBUS_OUT(121),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(121),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(121), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(122),
	GlitchData    => PPCMPLBWRDBUS122_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(122)",
	OutTemp       => PPCMPLBWRDBUS_OUT(122),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(122),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(122), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(123),
	GlitchData    => PPCMPLBWRDBUS123_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(123)",
	OutTemp       => PPCMPLBWRDBUS_OUT(123),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(123),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(123), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(124),
	GlitchData    => PPCMPLBWRDBUS124_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(124)",
	OutTemp       => PPCMPLBWRDBUS_OUT(124),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(124),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(124), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(125),
	GlitchData    => PPCMPLBWRDBUS125_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(125)",
	OutTemp       => PPCMPLBWRDBUS_OUT(125),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(125),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(125), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(126),
	GlitchData    => PPCMPLBWRDBUS126_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(126)",
	OutTemp       => PPCMPLBWRDBUS_OUT(126),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(126),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(126), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCMPLBWRDBUS(127),
	GlitchData    => PPCMPLBWRDBUS127_GlitchData,
	OutSignalName => "PPCMPLBWRDBUS(127)",
	OutTemp       => PPCMPLBWRDBUS_OUT(127),
	Paths       => (0 => (CPMPPCMPLBCLK_dly'last_event, tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(127),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCMPLBCLK_PPCMPLBWRDBUS(127), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBADDRACK,
	GlitchData    => PPCS0PLBADDRACK_GlitchData,
	OutSignalName => "PPCS0PLBADDRACK",
	OutTemp       => PPCS0PLBADDRACK_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBADDRACK,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBADDRACK, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMBUSY(0),
	GlitchData    => PPCS0PLBMBUSY0_GlitchData,
	OutSignalName => "PPCS0PLBMBUSY(0)",
	OutTemp       => PPCS0PLBMBUSY_OUT(0),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMBUSY(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMBUSY(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMBUSY(1),
	GlitchData    => PPCS0PLBMBUSY1_GlitchData,
	OutSignalName => "PPCS0PLBMBUSY(1)",
	OutTemp       => PPCS0PLBMBUSY_OUT(1),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMBUSY(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMBUSY(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMBUSY(2),
	GlitchData    => PPCS0PLBMBUSY2_GlitchData,
	OutSignalName => "PPCS0PLBMBUSY(2)",
	OutTemp       => PPCS0PLBMBUSY_OUT(2),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMBUSY(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMBUSY(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMBUSY(3),
	GlitchData    => PPCS0PLBMBUSY3_GlitchData,
	OutSignalName => "PPCS0PLBMBUSY(3)",
	OutTemp       => PPCS0PLBMBUSY_OUT(3),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMBUSY(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMBUSY(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMIRQ(0),
	GlitchData    => PPCS0PLBMIRQ0_GlitchData,
	OutSignalName => "PPCS0PLBMIRQ(0)",
	OutTemp       => PPCS0PLBMIRQ_OUT(0),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMIRQ(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMIRQ(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMIRQ(1),
	GlitchData    => PPCS0PLBMIRQ1_GlitchData,
	OutSignalName => "PPCS0PLBMIRQ(1)",
	OutTemp       => PPCS0PLBMIRQ_OUT(1),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMIRQ(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMIRQ(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMIRQ(2),
	GlitchData    => PPCS0PLBMIRQ2_GlitchData,
	OutSignalName => "PPCS0PLBMIRQ(2)",
	OutTemp       => PPCS0PLBMIRQ_OUT(2),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMIRQ(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMIRQ(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMIRQ(3),
	GlitchData    => PPCS0PLBMIRQ3_GlitchData,
	OutSignalName => "PPCS0PLBMIRQ(3)",
	OutTemp       => PPCS0PLBMIRQ_OUT(3),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMIRQ(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMIRQ(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMRDERR(0),
	GlitchData    => PPCS0PLBMRDERR0_GlitchData,
	OutSignalName => "PPCS0PLBMRDERR(0)",
	OutTemp       => PPCS0PLBMRDERR_OUT(0),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMRDERR(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMRDERR(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMRDERR(1),
	GlitchData    => PPCS0PLBMRDERR1_GlitchData,
	OutSignalName => "PPCS0PLBMRDERR(1)",
	OutTemp       => PPCS0PLBMRDERR_OUT(1),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMRDERR(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMRDERR(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMRDERR(2),
	GlitchData    => PPCS0PLBMRDERR2_GlitchData,
	OutSignalName => "PPCS0PLBMRDERR(2)",
	OutTemp       => PPCS0PLBMRDERR_OUT(2),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMRDERR(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMRDERR(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMRDERR(3),
	GlitchData    => PPCS0PLBMRDERR3_GlitchData,
	OutSignalName => "PPCS0PLBMRDERR(3)",
	OutTemp       => PPCS0PLBMRDERR_OUT(3),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMRDERR(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMRDERR(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMWRERR(0),
	GlitchData    => PPCS0PLBMWRERR0_GlitchData,
	OutSignalName => "PPCS0PLBMWRERR(0)",
	OutTemp       => PPCS0PLBMWRERR_OUT(0),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMWRERR(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMWRERR(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMWRERR(1),
	GlitchData    => PPCS0PLBMWRERR1_GlitchData,
	OutSignalName => "PPCS0PLBMWRERR(1)",
	OutTemp       => PPCS0PLBMWRERR_OUT(1),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMWRERR(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMWRERR(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMWRERR(2),
	GlitchData    => PPCS0PLBMWRERR2_GlitchData,
	OutSignalName => "PPCS0PLBMWRERR(2)",
	OutTemp       => PPCS0PLBMWRERR_OUT(2),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMWRERR(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMWRERR(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBMWRERR(3),
	GlitchData    => PPCS0PLBMWRERR3_GlitchData,
	OutSignalName => "PPCS0PLBMWRERR(3)",
	OutTemp       => PPCS0PLBMWRERR_OUT(3),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBMWRERR(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBMWRERR(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDBTERM,
	GlitchData    => PPCS0PLBRDBTERM_GlitchData,
	OutSignalName => "PPCS0PLBRDBTERM",
	OutTemp       => PPCS0PLBRDBTERM_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDBTERM,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDBTERM, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDCOMP,
	GlitchData    => PPCS0PLBRDCOMP_GlitchData,
	OutSignalName => "PPCS0PLBRDCOMP",
	OutTemp       => PPCS0PLBRDCOMP_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDCOMP,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDCOMP, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDACK,
	GlitchData    => PPCS0PLBRDDACK_GlitchData,
	OutSignalName => "PPCS0PLBRDDACK",
	OutTemp       => PPCS0PLBRDDACK_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDACK,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDACK, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(0),
	GlitchData    => PPCS0PLBRDDBUS0_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(0)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(0),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(1),
	GlitchData    => PPCS0PLBRDDBUS1_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(1)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(1),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(2),
	GlitchData    => PPCS0PLBRDDBUS2_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(2)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(2),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(3),
	GlitchData    => PPCS0PLBRDDBUS3_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(3)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(3),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(4),
	GlitchData    => PPCS0PLBRDDBUS4_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(4)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(4),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(4),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(5),
	GlitchData    => PPCS0PLBRDDBUS5_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(5)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(5),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(5),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(6),
	GlitchData    => PPCS0PLBRDDBUS6_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(6)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(6),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(6),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(7),
	GlitchData    => PPCS0PLBRDDBUS7_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(7)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(7),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(7),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(8),
	GlitchData    => PPCS0PLBRDDBUS8_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(8)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(8),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(8),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(9),
	GlitchData    => PPCS0PLBRDDBUS9_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(9)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(9),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(9),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(10),
	GlitchData    => PPCS0PLBRDDBUS10_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(10)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(10),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(10),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(11),
	GlitchData    => PPCS0PLBRDDBUS11_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(11)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(11),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(11),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(12),
	GlitchData    => PPCS0PLBRDDBUS12_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(12)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(12),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(12),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(13),
	GlitchData    => PPCS0PLBRDDBUS13_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(13)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(13),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(13),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(14),
	GlitchData    => PPCS0PLBRDDBUS14_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(14)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(14),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(14),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(15),
	GlitchData    => PPCS0PLBRDDBUS15_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(15)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(15),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(15),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(16),
	GlitchData    => PPCS0PLBRDDBUS16_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(16)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(16),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(16),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(17),
	GlitchData    => PPCS0PLBRDDBUS17_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(17)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(17),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(17),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(18),
	GlitchData    => PPCS0PLBRDDBUS18_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(18)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(18),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(18),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(19),
	GlitchData    => PPCS0PLBRDDBUS19_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(19)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(19),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(19),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(20),
	GlitchData    => PPCS0PLBRDDBUS20_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(20)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(20),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(20),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(21),
	GlitchData    => PPCS0PLBRDDBUS21_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(21)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(21),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(21),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(22),
	GlitchData    => PPCS0PLBRDDBUS22_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(22)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(22),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(22),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(23),
	GlitchData    => PPCS0PLBRDDBUS23_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(23)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(23),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(23),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(24),
	GlitchData    => PPCS0PLBRDDBUS24_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(24)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(24),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(24),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(25),
	GlitchData    => PPCS0PLBRDDBUS25_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(25)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(25),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(25),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(26),
	GlitchData    => PPCS0PLBRDDBUS26_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(26)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(26),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(26),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(27),
	GlitchData    => PPCS0PLBRDDBUS27_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(27)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(27),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(27),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(28),
	GlitchData    => PPCS0PLBRDDBUS28_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(28)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(28),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(28),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(29),
	GlitchData    => PPCS0PLBRDDBUS29_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(29)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(29),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(29),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(30),
	GlitchData    => PPCS0PLBRDDBUS30_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(30)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(30),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(30),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(31),
	GlitchData    => PPCS0PLBRDDBUS31_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(31)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(31),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(31),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(32),
	GlitchData    => PPCS0PLBRDDBUS32_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(32)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(32),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(32),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(32), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(33),
	GlitchData    => PPCS0PLBRDDBUS33_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(33)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(33),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(33),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(33), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(34),
	GlitchData    => PPCS0PLBRDDBUS34_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(34)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(34),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(34),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(34), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(35),
	GlitchData    => PPCS0PLBRDDBUS35_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(35)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(35),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(35),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(35), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(36),
	GlitchData    => PPCS0PLBRDDBUS36_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(36)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(36),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(36),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(36), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(37),
	GlitchData    => PPCS0PLBRDDBUS37_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(37)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(37),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(37),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(37), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(38),
	GlitchData    => PPCS0PLBRDDBUS38_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(38)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(38),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(38),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(38), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(39),
	GlitchData    => PPCS0PLBRDDBUS39_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(39)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(39),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(39),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(39), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(40),
	GlitchData    => PPCS0PLBRDDBUS40_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(40)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(40),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(40),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(40), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(41),
	GlitchData    => PPCS0PLBRDDBUS41_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(41)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(41),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(41),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(41), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(42),
	GlitchData    => PPCS0PLBRDDBUS42_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(42)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(42),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(42),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(42), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(43),
	GlitchData    => PPCS0PLBRDDBUS43_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(43)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(43),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(43),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(43), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(44),
	GlitchData    => PPCS0PLBRDDBUS44_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(44)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(44),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(44),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(44), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(45),
	GlitchData    => PPCS0PLBRDDBUS45_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(45)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(45),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(45),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(45), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(46),
	GlitchData    => PPCS0PLBRDDBUS46_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(46)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(46),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(46),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(46), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(47),
	GlitchData    => PPCS0PLBRDDBUS47_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(47)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(47),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(47),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(47), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(48),
	GlitchData    => PPCS0PLBRDDBUS48_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(48)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(48),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(48),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(48), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(49),
	GlitchData    => PPCS0PLBRDDBUS49_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(49)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(49),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(49),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(49), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(50),
	GlitchData    => PPCS0PLBRDDBUS50_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(50)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(50),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(50),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(50), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(51),
	GlitchData    => PPCS0PLBRDDBUS51_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(51)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(51),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(51),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(51), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(52),
	GlitchData    => PPCS0PLBRDDBUS52_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(52)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(52),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(52),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(52), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(53),
	GlitchData    => PPCS0PLBRDDBUS53_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(53)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(53),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(53),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(53), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(54),
	GlitchData    => PPCS0PLBRDDBUS54_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(54)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(54),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(54),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(54), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(55),
	GlitchData    => PPCS0PLBRDDBUS55_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(55)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(55),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(55),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(55), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(56),
	GlitchData    => PPCS0PLBRDDBUS56_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(56)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(56),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(56),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(56), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(57),
	GlitchData    => PPCS0PLBRDDBUS57_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(57)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(57),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(57),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(57), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(58),
	GlitchData    => PPCS0PLBRDDBUS58_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(58)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(58),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(58),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(58), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(59),
	GlitchData    => PPCS0PLBRDDBUS59_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(59)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(59),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(59),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(59), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(60),
	GlitchData    => PPCS0PLBRDDBUS60_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(60)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(60),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(60),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(60), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(61),
	GlitchData    => PPCS0PLBRDDBUS61_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(61)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(61),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(61),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(61), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(62),
	GlitchData    => PPCS0PLBRDDBUS62_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(62)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(62),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(62),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(62), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(63),
	GlitchData    => PPCS0PLBRDDBUS63_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(63)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(63),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(63),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(63), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(64),
	GlitchData    => PPCS0PLBRDDBUS64_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(64)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(64),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(64),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(64), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(65),
	GlitchData    => PPCS0PLBRDDBUS65_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(65)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(65),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(65),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(65), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(66),
	GlitchData    => PPCS0PLBRDDBUS66_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(66)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(66),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(66),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(66), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(67),
	GlitchData    => PPCS0PLBRDDBUS67_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(67)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(67),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(67),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(67), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(68),
	GlitchData    => PPCS0PLBRDDBUS68_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(68)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(68),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(68),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(68), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(69),
	GlitchData    => PPCS0PLBRDDBUS69_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(69)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(69),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(69),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(69), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(70),
	GlitchData    => PPCS0PLBRDDBUS70_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(70)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(70),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(70),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(70), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(71),
	GlitchData    => PPCS0PLBRDDBUS71_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(71)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(71),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(71),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(71), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(72),
	GlitchData    => PPCS0PLBRDDBUS72_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(72)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(72),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(72),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(72), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(73),
	GlitchData    => PPCS0PLBRDDBUS73_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(73)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(73),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(73),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(73), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(74),
	GlitchData    => PPCS0PLBRDDBUS74_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(74)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(74),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(74),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(74), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(75),
	GlitchData    => PPCS0PLBRDDBUS75_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(75)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(75),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(75),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(75), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(76),
	GlitchData    => PPCS0PLBRDDBUS76_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(76)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(76),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(76),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(76), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(77),
	GlitchData    => PPCS0PLBRDDBUS77_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(77)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(77),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(77),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(77), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(78),
	GlitchData    => PPCS0PLBRDDBUS78_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(78)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(78),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(78),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(78), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(79),
	GlitchData    => PPCS0PLBRDDBUS79_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(79)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(79),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(79),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(79), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(80),
	GlitchData    => PPCS0PLBRDDBUS80_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(80)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(80),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(80),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(80), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(81),
	GlitchData    => PPCS0PLBRDDBUS81_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(81)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(81),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(81),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(81), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(82),
	GlitchData    => PPCS0PLBRDDBUS82_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(82)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(82),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(82),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(82), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(83),
	GlitchData    => PPCS0PLBRDDBUS83_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(83)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(83),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(83),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(83), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(84),
	GlitchData    => PPCS0PLBRDDBUS84_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(84)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(84),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(84),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(84), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(85),
	GlitchData    => PPCS0PLBRDDBUS85_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(85)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(85),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(85),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(85), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(86),
	GlitchData    => PPCS0PLBRDDBUS86_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(86)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(86),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(86),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(86), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(87),
	GlitchData    => PPCS0PLBRDDBUS87_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(87)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(87),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(87),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(87), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(88),
	GlitchData    => PPCS0PLBRDDBUS88_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(88)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(88),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(88),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(88), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(89),
	GlitchData    => PPCS0PLBRDDBUS89_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(89)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(89),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(89),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(89), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(90),
	GlitchData    => PPCS0PLBRDDBUS90_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(90)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(90),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(90),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(90), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(91),
	GlitchData    => PPCS0PLBRDDBUS91_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(91)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(91),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(91),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(91), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(92),
	GlitchData    => PPCS0PLBRDDBUS92_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(92)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(92),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(92),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(92), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(93),
	GlitchData    => PPCS0PLBRDDBUS93_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(93)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(93),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(93),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(93), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(94),
	GlitchData    => PPCS0PLBRDDBUS94_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(94)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(94),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(94),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(94), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(95),
	GlitchData    => PPCS0PLBRDDBUS95_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(95)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(95),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(95),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(95), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(96),
	GlitchData    => PPCS0PLBRDDBUS96_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(96)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(96),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(96),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(96), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(97),
	GlitchData    => PPCS0PLBRDDBUS97_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(97)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(97),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(97),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(97), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(98),
	GlitchData    => PPCS0PLBRDDBUS98_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(98)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(98),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(98),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(98), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(99),
	GlitchData    => PPCS0PLBRDDBUS99_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(99)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(99),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(99),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(99), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(100),
	GlitchData    => PPCS0PLBRDDBUS100_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(100)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(100),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(100),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(100), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(101),
	GlitchData    => PPCS0PLBRDDBUS101_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(101)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(101),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(101),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(101), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(102),
	GlitchData    => PPCS0PLBRDDBUS102_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(102)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(102),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(102),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(102), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(103),
	GlitchData    => PPCS0PLBRDDBUS103_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(103)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(103),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(103),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(103), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(104),
	GlitchData    => PPCS0PLBRDDBUS104_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(104)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(104),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(104),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(104), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(105),
	GlitchData    => PPCS0PLBRDDBUS105_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(105)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(105),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(105),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(105), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(106),
	GlitchData    => PPCS0PLBRDDBUS106_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(106)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(106),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(106),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(106), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(107),
	GlitchData    => PPCS0PLBRDDBUS107_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(107)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(107),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(107),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(107), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(108),
	GlitchData    => PPCS0PLBRDDBUS108_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(108)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(108),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(108),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(108), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(109),
	GlitchData    => PPCS0PLBRDDBUS109_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(109)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(109),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(109),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(109), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(110),
	GlitchData    => PPCS0PLBRDDBUS110_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(110)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(110),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(110),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(110), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(111),
	GlitchData    => PPCS0PLBRDDBUS111_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(111)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(111),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(111),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(111), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(112),
	GlitchData    => PPCS0PLBRDDBUS112_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(112)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(112),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(112),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(112), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(113),
	GlitchData    => PPCS0PLBRDDBUS113_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(113)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(113),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(113),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(113), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(114),
	GlitchData    => PPCS0PLBRDDBUS114_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(114)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(114),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(114),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(114), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(115),
	GlitchData    => PPCS0PLBRDDBUS115_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(115)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(115),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(115),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(115), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(116),
	GlitchData    => PPCS0PLBRDDBUS116_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(116)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(116),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(116),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(116), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(117),
	GlitchData    => PPCS0PLBRDDBUS117_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(117)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(117),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(117),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(117), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(118),
	GlitchData    => PPCS0PLBRDDBUS118_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(118)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(118),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(118),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(118), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(119),
	GlitchData    => PPCS0PLBRDDBUS119_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(119)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(119),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(119),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(119), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(120),
	GlitchData    => PPCS0PLBRDDBUS120_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(120)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(120),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(120),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(120), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(121),
	GlitchData    => PPCS0PLBRDDBUS121_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(121)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(121),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(121),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(121), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(122),
	GlitchData    => PPCS0PLBRDDBUS122_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(122)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(122),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(122),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(122), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(123),
	GlitchData    => PPCS0PLBRDDBUS123_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(123)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(123),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(123),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(123), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(124),
	GlitchData    => PPCS0PLBRDDBUS124_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(124)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(124),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(124),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(124), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(125),
	GlitchData    => PPCS0PLBRDDBUS125_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(125)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(125),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(125),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(125), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(126),
	GlitchData    => PPCS0PLBRDDBUS126_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(126)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(126),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(126),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(126), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDDBUS(127),
	GlitchData    => PPCS0PLBRDDBUS127_GlitchData,
	OutSignalName => "PPCS0PLBRDDBUS(127)",
	OutTemp       => PPCS0PLBRDDBUS_OUT(127),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(127),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDDBUS(127), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDWDADDR(0),
	GlitchData    => PPCS0PLBRDWDADDR0_GlitchData,
	OutSignalName => "PPCS0PLBRDWDADDR(0)",
	OutTemp       => PPCS0PLBRDWDADDR_OUT(0),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDWDADDR(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDWDADDR(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDWDADDR(1),
	GlitchData    => PPCS0PLBRDWDADDR1_GlitchData,
	OutSignalName => "PPCS0PLBRDWDADDR(1)",
	OutTemp       => PPCS0PLBRDWDADDR_OUT(1),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDWDADDR(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDWDADDR(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDWDADDR(2),
	GlitchData    => PPCS0PLBRDWDADDR2_GlitchData,
	OutSignalName => "PPCS0PLBRDWDADDR(2)",
	OutTemp       => PPCS0PLBRDWDADDR_OUT(2),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDWDADDR(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDWDADDR(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBRDWDADDR(3),
	GlitchData    => PPCS0PLBRDWDADDR3_GlitchData,
	OutSignalName => "PPCS0PLBRDWDADDR(3)",
	OutTemp       => PPCS0PLBRDWDADDR_OUT(3),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBRDWDADDR(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBRDWDADDR(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBREARBITRATE,
	GlitchData    => PPCS0PLBREARBITRATE_GlitchData,
	OutSignalName => "PPCS0PLBREARBITRATE",
	OutTemp       => PPCS0PLBREARBITRATE_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBREARBITRATE,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBREARBITRATE, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBSSIZE(0),
	GlitchData    => PPCS0PLBSSIZE0_GlitchData,
	OutSignalName => "PPCS0PLBSSIZE(0)",
	OutTemp       => PPCS0PLBSSIZE_OUT(0),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBSSIZE(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBSSIZE(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBSSIZE(1),
	GlitchData    => PPCS0PLBSSIZE1_GlitchData,
	OutSignalName => "PPCS0PLBSSIZE(1)",
	OutTemp       => PPCS0PLBSSIZE_OUT(1),
	Paths       => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBSSIZE(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBSSIZE(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBWAIT,
	GlitchData    => PPCS0PLBWAIT_GlitchData,
	OutSignalName => "PPCS0PLBWAIT",
	OutTemp       => PPCS0PLBWAIT_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBWAIT,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBWAIT, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBWRBTERM,
	GlitchData    => PPCS0PLBWRBTERM_GlitchData,
	OutSignalName => "PPCS0PLBWRBTERM",
	OutTemp       => PPCS0PLBWRBTERM_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBWRBTERM,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBWRBTERM, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBWRCOMP,
	GlitchData    => PPCS0PLBWRCOMP_GlitchData,
	OutSignalName => "PPCS0PLBWRCOMP",
	OutTemp       => PPCS0PLBWRCOMP_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBWRCOMP,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBWRCOMP, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS0PLBWRDACK,
	GlitchData    => PPCS0PLBWRDACK_GlitchData,
	OutSignalName => "PPCS0PLBWRDACK",
	OutTemp       => PPCS0PLBWRDACK_OUT,
	Paths         => (0 => (CPMPPCS0PLBCLK_dly'last_event, tpd_CPMPPCS0PLBCLK_PPCS0PLBWRDACK,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS0PLBCLK_PPCS0PLBWRDACK, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBADDRACK,
	GlitchData    => PPCS1PLBADDRACK_GlitchData,
	OutSignalName => "PPCS1PLBADDRACK",
	OutTemp       => PPCS1PLBADDRACK_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBADDRACK,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBADDRACK, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMBUSY(0),
	GlitchData    => PPCS1PLBMBUSY0_GlitchData,
	OutSignalName => "PPCS1PLBMBUSY(0)",
	OutTemp       => PPCS1PLBMBUSY_OUT(0),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMBUSY(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMBUSY(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMBUSY(1),
	GlitchData    => PPCS1PLBMBUSY1_GlitchData,
	OutSignalName => "PPCS1PLBMBUSY(1)",
	OutTemp       => PPCS1PLBMBUSY_OUT(1),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMBUSY(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMBUSY(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMBUSY(2),
	GlitchData    => PPCS1PLBMBUSY2_GlitchData,
	OutSignalName => "PPCS1PLBMBUSY(2)",
	OutTemp       => PPCS1PLBMBUSY_OUT(2),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMBUSY(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMBUSY(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMBUSY(3),
	GlitchData    => PPCS1PLBMBUSY3_GlitchData,
	OutSignalName => "PPCS1PLBMBUSY(3)",
	OutTemp       => PPCS1PLBMBUSY_OUT(3),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMBUSY(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMBUSY(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMIRQ(0),
	GlitchData    => PPCS1PLBMIRQ0_GlitchData,
	OutSignalName => "PPCS1PLBMIRQ(0)",
	OutTemp       => PPCS1PLBMIRQ_OUT(0),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMIRQ(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMIRQ(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMIRQ(1),
	GlitchData    => PPCS1PLBMIRQ1_GlitchData,
	OutSignalName => "PPCS1PLBMIRQ(1)",
	OutTemp       => PPCS1PLBMIRQ_OUT(1),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMIRQ(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMIRQ(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMIRQ(2),
	GlitchData    => PPCS1PLBMIRQ2_GlitchData,
	OutSignalName => "PPCS1PLBMIRQ(2)",
	OutTemp       => PPCS1PLBMIRQ_OUT(2),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMIRQ(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMIRQ(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMIRQ(3),
	GlitchData    => PPCS1PLBMIRQ3_GlitchData,
	OutSignalName => "PPCS1PLBMIRQ(3)",
	OutTemp       => PPCS1PLBMIRQ_OUT(3),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMIRQ(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMIRQ(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMRDERR(0),
	GlitchData    => PPCS1PLBMRDERR0_GlitchData,
	OutSignalName => "PPCS1PLBMRDERR(0)",
	OutTemp       => PPCS1PLBMRDERR_OUT(0),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMRDERR(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMRDERR(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMRDERR(1),
	GlitchData    => PPCS1PLBMRDERR1_GlitchData,
	OutSignalName => "PPCS1PLBMRDERR(1)",
	OutTemp       => PPCS1PLBMRDERR_OUT(1),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMRDERR(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMRDERR(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMRDERR(2),
	GlitchData    => PPCS1PLBMRDERR2_GlitchData,
	OutSignalName => "PPCS1PLBMRDERR(2)",
	OutTemp       => PPCS1PLBMRDERR_OUT(2),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMRDERR(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMRDERR(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMRDERR(3),
	GlitchData    => PPCS1PLBMRDERR3_GlitchData,
	OutSignalName => "PPCS1PLBMRDERR(3)",
	OutTemp       => PPCS1PLBMRDERR_OUT(3),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMRDERR(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMRDERR(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMWRERR(0),
	GlitchData    => PPCS1PLBMWRERR0_GlitchData,
	OutSignalName => "PPCS1PLBMWRERR(0)",
	OutTemp       => PPCS1PLBMWRERR_OUT(0),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMWRERR(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMWRERR(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMWRERR(1),
	GlitchData    => PPCS1PLBMWRERR1_GlitchData,
	OutSignalName => "PPCS1PLBMWRERR(1)",
	OutTemp       => PPCS1PLBMWRERR_OUT(1),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMWRERR(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMWRERR(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMWRERR(2),
	GlitchData    => PPCS1PLBMWRERR2_GlitchData,
	OutSignalName => "PPCS1PLBMWRERR(2)",
	OutTemp       => PPCS1PLBMWRERR_OUT(2),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMWRERR(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMWRERR(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBMWRERR(3),
	GlitchData    => PPCS1PLBMWRERR3_GlitchData,
	OutSignalName => "PPCS1PLBMWRERR(3)",
	OutTemp       => PPCS1PLBMWRERR_OUT(3),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBMWRERR(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBMWRERR(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDBTERM,
	GlitchData    => PPCS1PLBRDBTERM_GlitchData,
	OutSignalName => "PPCS1PLBRDBTERM",
	OutTemp       => PPCS1PLBRDBTERM_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDBTERM,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDBTERM, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDCOMP,
	GlitchData    => PPCS1PLBRDCOMP_GlitchData,
	OutSignalName => "PPCS1PLBRDCOMP",
	OutTemp       => PPCS1PLBRDCOMP_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDCOMP,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDCOMP, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDACK,
	GlitchData    => PPCS1PLBRDDACK_GlitchData,
	OutSignalName => "PPCS1PLBRDDACK",
	OutTemp       => PPCS1PLBRDDACK_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDACK,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDACK, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(0),
	GlitchData    => PPCS1PLBRDDBUS0_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(0)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(0),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(1),
	GlitchData    => PPCS1PLBRDDBUS1_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(1)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(1),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(2),
	GlitchData    => PPCS1PLBRDDBUS2_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(2)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(2),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(3),
	GlitchData    => PPCS1PLBRDDBUS3_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(3)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(3),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(4),
	GlitchData    => PPCS1PLBRDDBUS4_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(4)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(4),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(4),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(5),
	GlitchData    => PPCS1PLBRDDBUS5_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(5)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(5),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(5),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(6),
	GlitchData    => PPCS1PLBRDDBUS6_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(6)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(6),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(6),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(7),
	GlitchData    => PPCS1PLBRDDBUS7_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(7)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(7),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(7),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(8),
	GlitchData    => PPCS1PLBRDDBUS8_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(8)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(8),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(8),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(9),
	GlitchData    => PPCS1PLBRDDBUS9_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(9)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(9),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(9),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(10),
	GlitchData    => PPCS1PLBRDDBUS10_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(10)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(10),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(10),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(11),
	GlitchData    => PPCS1PLBRDDBUS11_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(11)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(11),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(11),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(12),
	GlitchData    => PPCS1PLBRDDBUS12_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(12)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(12),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(12),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(13),
	GlitchData    => PPCS1PLBRDDBUS13_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(13)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(13),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(13),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(14),
	GlitchData    => PPCS1PLBRDDBUS14_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(14)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(14),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(14),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(15),
	GlitchData    => PPCS1PLBRDDBUS15_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(15)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(15),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(15),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(16),
	GlitchData    => PPCS1PLBRDDBUS16_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(16)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(16),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(16),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(17),
	GlitchData    => PPCS1PLBRDDBUS17_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(17)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(17),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(17),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(18),
	GlitchData    => PPCS1PLBRDDBUS18_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(18)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(18),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(18),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(19),
	GlitchData    => PPCS1PLBRDDBUS19_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(19)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(19),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(19),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(20),
	GlitchData    => PPCS1PLBRDDBUS20_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(20)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(20),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(20),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(21),
	GlitchData    => PPCS1PLBRDDBUS21_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(21)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(21),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(21),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(22),
	GlitchData    => PPCS1PLBRDDBUS22_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(22)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(22),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(22),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(23),
	GlitchData    => PPCS1PLBRDDBUS23_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(23)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(23),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(23),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(24),
	GlitchData    => PPCS1PLBRDDBUS24_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(24)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(24),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(24),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(25),
	GlitchData    => PPCS1PLBRDDBUS25_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(25)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(25),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(25),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(26),
	GlitchData    => PPCS1PLBRDDBUS26_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(26)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(26),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(26),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(27),
	GlitchData    => PPCS1PLBRDDBUS27_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(27)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(27),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(27),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(28),
	GlitchData    => PPCS1PLBRDDBUS28_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(28)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(28),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(28),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(29),
	GlitchData    => PPCS1PLBRDDBUS29_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(29)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(29),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(29),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(30),
	GlitchData    => PPCS1PLBRDDBUS30_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(30)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(30),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(30),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(31),
	GlitchData    => PPCS1PLBRDDBUS31_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(31)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(31),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(31),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(32),
	GlitchData    => PPCS1PLBRDDBUS32_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(32)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(32),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(32),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(32), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(33),
	GlitchData    => PPCS1PLBRDDBUS33_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(33)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(33),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(33),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(33), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(34),
	GlitchData    => PPCS1PLBRDDBUS34_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(34)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(34),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(34),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(34), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(35),
	GlitchData    => PPCS1PLBRDDBUS35_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(35)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(35),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(35),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(35), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(36),
	GlitchData    => PPCS1PLBRDDBUS36_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(36)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(36),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(36),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(36), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(37),
	GlitchData    => PPCS1PLBRDDBUS37_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(37)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(37),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(37),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(37), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(38),
	GlitchData    => PPCS1PLBRDDBUS38_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(38)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(38),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(38),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(38), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(39),
	GlitchData    => PPCS1PLBRDDBUS39_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(39)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(39),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(39),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(39), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(40),
	GlitchData    => PPCS1PLBRDDBUS40_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(40)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(40),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(40),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(40), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(41),
	GlitchData    => PPCS1PLBRDDBUS41_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(41)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(41),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(41),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(41), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(42),
	GlitchData    => PPCS1PLBRDDBUS42_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(42)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(42),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(42),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(42), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(43),
	GlitchData    => PPCS1PLBRDDBUS43_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(43)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(43),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(43),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(43), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(44),
	GlitchData    => PPCS1PLBRDDBUS44_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(44)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(44),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(44),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(44), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(45),
	GlitchData    => PPCS1PLBRDDBUS45_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(45)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(45),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(45),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(45), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(46),
	GlitchData    => PPCS1PLBRDDBUS46_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(46)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(46),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(46),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(46), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(47),
	GlitchData    => PPCS1PLBRDDBUS47_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(47)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(47),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(47),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(47), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(48),
	GlitchData    => PPCS1PLBRDDBUS48_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(48)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(48),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(48),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(48), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(49),
	GlitchData    => PPCS1PLBRDDBUS49_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(49)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(49),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(49),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(49), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(50),
	GlitchData    => PPCS1PLBRDDBUS50_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(50)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(50),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(50),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(50), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(51),
	GlitchData    => PPCS1PLBRDDBUS51_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(51)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(51),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(51),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(51), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(52),
	GlitchData    => PPCS1PLBRDDBUS52_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(52)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(52),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(52),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(52), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(53),
	GlitchData    => PPCS1PLBRDDBUS53_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(53)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(53),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(53),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(53), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(54),
	GlitchData    => PPCS1PLBRDDBUS54_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(54)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(54),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(54),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(54), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(55),
	GlitchData    => PPCS1PLBRDDBUS55_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(55)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(55),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(55),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(55), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(56),
	GlitchData    => PPCS1PLBRDDBUS56_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(56)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(56),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(56),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(56), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(57),
	GlitchData    => PPCS1PLBRDDBUS57_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(57)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(57),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(57),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(57), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(58),
	GlitchData    => PPCS1PLBRDDBUS58_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(58)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(58),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(58),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(58), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(59),
	GlitchData    => PPCS1PLBRDDBUS59_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(59)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(59),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(59),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(59), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(60),
	GlitchData    => PPCS1PLBRDDBUS60_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(60)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(60),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(60),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(60), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(61),
	GlitchData    => PPCS1PLBRDDBUS61_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(61)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(61),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(61),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(61), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(62),
	GlitchData    => PPCS1PLBRDDBUS62_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(62)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(62),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(62),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(62), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(63),
	GlitchData    => PPCS1PLBRDDBUS63_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(63)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(63),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(63),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(63), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(64),
	GlitchData    => PPCS1PLBRDDBUS64_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(64)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(64),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(64),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(64), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(65),
	GlitchData    => PPCS1PLBRDDBUS65_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(65)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(65),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(65),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(65), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(66),
	GlitchData    => PPCS1PLBRDDBUS66_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(66)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(66),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(66),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(66), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(67),
	GlitchData    => PPCS1PLBRDDBUS67_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(67)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(67),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(67),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(67), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(68),
	GlitchData    => PPCS1PLBRDDBUS68_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(68)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(68),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(68),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(68), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(69),
	GlitchData    => PPCS1PLBRDDBUS69_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(69)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(69),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(69),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(69), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(70),
	GlitchData    => PPCS1PLBRDDBUS70_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(70)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(70),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(70),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(70), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(71),
	GlitchData    => PPCS1PLBRDDBUS71_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(71)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(71),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(71),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(71), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(72),
	GlitchData    => PPCS1PLBRDDBUS72_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(72)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(72),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(72),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(72), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(73),
	GlitchData    => PPCS1PLBRDDBUS73_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(73)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(73),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(73),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(73), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(74),
	GlitchData    => PPCS1PLBRDDBUS74_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(74)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(74),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(74),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(74), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(75),
	GlitchData    => PPCS1PLBRDDBUS75_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(75)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(75),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(75),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(75), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(76),
	GlitchData    => PPCS1PLBRDDBUS76_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(76)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(76),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(76),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(76), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(77),
	GlitchData    => PPCS1PLBRDDBUS77_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(77)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(77),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(77),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(77), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(78),
	GlitchData    => PPCS1PLBRDDBUS78_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(78)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(78),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(78),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(78), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(79),
	GlitchData    => PPCS1PLBRDDBUS79_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(79)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(79),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(79),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(79), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(80),
	GlitchData    => PPCS1PLBRDDBUS80_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(80)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(80),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(80),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(80), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(81),
	GlitchData    => PPCS1PLBRDDBUS81_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(81)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(81),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(81),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(81), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(82),
	GlitchData    => PPCS1PLBRDDBUS82_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(82)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(82),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(82),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(82), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(83),
	GlitchData    => PPCS1PLBRDDBUS83_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(83)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(83),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(83),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(83), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(84),
	GlitchData    => PPCS1PLBRDDBUS84_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(84)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(84),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(84),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(84), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(85),
	GlitchData    => PPCS1PLBRDDBUS85_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(85)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(85),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(85),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(85), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(86),
	GlitchData    => PPCS1PLBRDDBUS86_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(86)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(86),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(86),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(86), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(87),
	GlitchData    => PPCS1PLBRDDBUS87_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(87)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(87),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(87),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(87), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(88),
	GlitchData    => PPCS1PLBRDDBUS88_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(88)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(88),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(88),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(88), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(89),
	GlitchData    => PPCS1PLBRDDBUS89_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(89)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(89),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(89),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(89), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(90),
	GlitchData    => PPCS1PLBRDDBUS90_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(90)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(90),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(90),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(90), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(91),
	GlitchData    => PPCS1PLBRDDBUS91_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(91)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(91),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(91),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(91), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(92),
	GlitchData    => PPCS1PLBRDDBUS92_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(92)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(92),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(92),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(92), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(93),
	GlitchData    => PPCS1PLBRDDBUS93_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(93)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(93),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(93),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(93), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(94),
	GlitchData    => PPCS1PLBRDDBUS94_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(94)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(94),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(94),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(94), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(95),
	GlitchData    => PPCS1PLBRDDBUS95_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(95)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(95),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(95),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(95), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(96),
	GlitchData    => PPCS1PLBRDDBUS96_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(96)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(96),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(96),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(96), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(97),
	GlitchData    => PPCS1PLBRDDBUS97_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(97)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(97),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(97),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(97), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(98),
	GlitchData    => PPCS1PLBRDDBUS98_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(98)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(98),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(98),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(98), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(99),
	GlitchData    => PPCS1PLBRDDBUS99_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(99)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(99),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(99),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(99), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(100),
	GlitchData    => PPCS1PLBRDDBUS100_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(100)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(100),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(100),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(100), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(101),
	GlitchData    => PPCS1PLBRDDBUS101_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(101)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(101),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(101),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(101), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(102),
	GlitchData    => PPCS1PLBRDDBUS102_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(102)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(102),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(102),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(102), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(103),
	GlitchData    => PPCS1PLBRDDBUS103_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(103)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(103),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(103),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(103), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(104),
	GlitchData    => PPCS1PLBRDDBUS104_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(104)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(104),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(104),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(104), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(105),
	GlitchData    => PPCS1PLBRDDBUS105_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(105)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(105),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(105),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(105), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(106),
	GlitchData    => PPCS1PLBRDDBUS106_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(106)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(106),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(106),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(106), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(107),
	GlitchData    => PPCS1PLBRDDBUS107_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(107)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(107),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(107),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(107), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(108),
	GlitchData    => PPCS1PLBRDDBUS108_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(108)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(108),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(108),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(108), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(109),
	GlitchData    => PPCS1PLBRDDBUS109_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(109)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(109),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(109),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(109), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(110),
	GlitchData    => PPCS1PLBRDDBUS110_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(110)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(110),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(110),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(110), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(111),
	GlitchData    => PPCS1PLBRDDBUS111_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(111)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(111),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(111),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(111), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(112),
	GlitchData    => PPCS1PLBRDDBUS112_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(112)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(112),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(112),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(112), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(113),
	GlitchData    => PPCS1PLBRDDBUS113_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(113)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(113),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(113),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(113), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(114),
	GlitchData    => PPCS1PLBRDDBUS114_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(114)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(114),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(114),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(114), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(115),
	GlitchData    => PPCS1PLBRDDBUS115_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(115)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(115),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(115),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(115), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(116),
	GlitchData    => PPCS1PLBRDDBUS116_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(116)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(116),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(116),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(116), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(117),
	GlitchData    => PPCS1PLBRDDBUS117_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(117)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(117),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(117),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(117), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(118),
	GlitchData    => PPCS1PLBRDDBUS118_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(118)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(118),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(118),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(118), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(119),
	GlitchData    => PPCS1PLBRDDBUS119_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(119)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(119),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(119),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(119), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(120),
	GlitchData    => PPCS1PLBRDDBUS120_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(120)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(120),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(120),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(120), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(121),
	GlitchData    => PPCS1PLBRDDBUS121_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(121)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(121),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(121),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(121), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(122),
	GlitchData    => PPCS1PLBRDDBUS122_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(122)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(122),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(122),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(122), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(123),
	GlitchData    => PPCS1PLBRDDBUS123_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(123)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(123),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(123),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(123), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(124),
	GlitchData    => PPCS1PLBRDDBUS124_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(124)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(124),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(124),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(124), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(125),
	GlitchData    => PPCS1PLBRDDBUS125_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(125)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(125),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(125),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(125), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(126),
	GlitchData    => PPCS1PLBRDDBUS126_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(126)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(126),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(126),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(126), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDDBUS(127),
	GlitchData    => PPCS1PLBRDDBUS127_GlitchData,
	OutSignalName => "PPCS1PLBRDDBUS(127)",
	OutTemp       => PPCS1PLBRDDBUS_OUT(127),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(127),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDDBUS(127), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDWDADDR(0),
	GlitchData    => PPCS1PLBRDWDADDR0_GlitchData,
	OutSignalName => "PPCS1PLBRDWDADDR(0)",
	OutTemp       => PPCS1PLBRDWDADDR_OUT(0),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDWDADDR(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDWDADDR(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDWDADDR(1),
	GlitchData    => PPCS1PLBRDWDADDR1_GlitchData,
	OutSignalName => "PPCS1PLBRDWDADDR(1)",
	OutTemp       => PPCS1PLBRDWDADDR_OUT(1),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDWDADDR(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDWDADDR(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDWDADDR(2),
	GlitchData    => PPCS1PLBRDWDADDR2_GlitchData,
	OutSignalName => "PPCS1PLBRDWDADDR(2)",
	OutTemp       => PPCS1PLBRDWDADDR_OUT(2),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDWDADDR(2),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDWDADDR(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBRDWDADDR(3),
	GlitchData    => PPCS1PLBRDWDADDR3_GlitchData,
	OutSignalName => "PPCS1PLBRDWDADDR(3)",
	OutTemp       => PPCS1PLBRDWDADDR_OUT(3),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBRDWDADDR(3),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBRDWDADDR(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBREARBITRATE,
	GlitchData    => PPCS1PLBREARBITRATE_GlitchData,
	OutSignalName => "PPCS1PLBREARBITRATE",
	OutTemp       => PPCS1PLBREARBITRATE_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBREARBITRATE,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBREARBITRATE, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBSSIZE(0),
	GlitchData    => PPCS1PLBSSIZE0_GlitchData,
	OutSignalName => "PPCS1PLBSSIZE(0)",
	OutTemp       => PPCS1PLBSSIZE_OUT(0),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBSSIZE(0),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBSSIZE(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBSSIZE(1),
	GlitchData    => PPCS1PLBSSIZE1_GlitchData,
	OutSignalName => "PPCS1PLBSSIZE(1)",
	OutTemp       => PPCS1PLBSSIZE_OUT(1),
	Paths       => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBSSIZE(1),TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBSSIZE(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBWAIT,
	GlitchData    => PPCS1PLBWAIT_GlitchData,
	OutSignalName => "PPCS1PLBWAIT",
	OutTemp       => PPCS1PLBWAIT_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBWAIT,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBWAIT, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBWRBTERM,
	GlitchData    => PPCS1PLBWRBTERM_GlitchData,
	OutSignalName => "PPCS1PLBWRBTERM",
	OutTemp       => PPCS1PLBWRBTERM_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBWRBTERM,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBWRBTERM, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBWRCOMP,
	GlitchData    => PPCS1PLBWRCOMP_GlitchData,
	OutSignalName => "PPCS1PLBWRCOMP",
	OutTemp       => PPCS1PLBWRCOMP_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBWRCOMP,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBWRCOMP, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCS1PLBWRDACK,
	GlitchData    => PPCS1PLBWRDACK_GlitchData,
	OutSignalName => "PPCS1PLBWRDACK",
	OutTemp       => PPCS1PLBWRDACK_OUT,
	Paths         => (0 => (CPMPPCS1PLBCLK_dly'last_event, tpd_CPMPPCS1PLBCLK_PPCS1PLBWRDACK,TRUE)),
	 DefaultDelay =>  tpd_CPMPPCS1PLBCLK_PPCS1PLBWRDACK, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECFPUOP,
	GlitchData    => APUFCMDECFPUOP_GlitchData,
	OutSignalName => "APUFCMDECFPUOP",
	OutTemp       => APUFCMDECFPUOP_OUT,
	Paths         => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMDECFPUOP,TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMDECFPUOP, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECLDSTXFERSIZE(0),
	GlitchData    => APUFCMDECLDSTXFERSIZE0_GlitchData,
	OutSignalName => "APUFCMDECLDSTXFERSIZE(0)",
	OutTemp       => APUFCMDECLDSTXFERSIZE_OUT(0),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMDECLDSTXFERSIZE(0),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMDECLDSTXFERSIZE(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECLDSTXFERSIZE(1),
	GlitchData    => APUFCMDECLDSTXFERSIZE1_GlitchData,
	OutSignalName => "APUFCMDECLDSTXFERSIZE(1)",
	OutTemp       => APUFCMDECLDSTXFERSIZE_OUT(1),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMDECLDSTXFERSIZE(1),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMDECLDSTXFERSIZE(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECLDSTXFERSIZE(2),
	GlitchData    => APUFCMDECLDSTXFERSIZE2_GlitchData,
	OutSignalName => "APUFCMDECLDSTXFERSIZE(2)",
	OutTemp       => APUFCMDECLDSTXFERSIZE_OUT(2),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMDECLDSTXFERSIZE(2),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMDECLDSTXFERSIZE(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECLOAD,
	GlitchData    => APUFCMDECLOAD_GlitchData,
	OutSignalName => "APUFCMDECLOAD",
	OutTemp       => APUFCMDECLOAD_OUT,
	Paths         => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMDECLOAD,TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMDECLOAD, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECNONAUTON,
	GlitchData    => APUFCMDECNONAUTON_GlitchData,
	OutSignalName => "APUFCMDECNONAUTON",
	OutTemp       => APUFCMDECNONAUTON_OUT,
	Paths         => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMDECNONAUTON,TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMDECNONAUTON, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECSTORE,
	GlitchData    => APUFCMDECSTORE_GlitchData,
	OutSignalName => "APUFCMDECSTORE",
	OutTemp       => APUFCMDECSTORE_OUT,
	Paths         => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMDECSTORE,TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMDECSTORE, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECUDI(0),
	GlitchData    => APUFCMDECUDI0_GlitchData,
	OutSignalName => "APUFCMDECUDI(0)",
	OutTemp       => APUFCMDECUDI_OUT(0),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMDECUDI(0),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMDECUDI(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECUDI(1),
	GlitchData    => APUFCMDECUDI1_GlitchData,
	OutSignalName => "APUFCMDECUDI(1)",
	OutTemp       => APUFCMDECUDI_OUT(1),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMDECUDI(1),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMDECUDI(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECUDI(2),
	GlitchData    => APUFCMDECUDI2_GlitchData,
	OutSignalName => "APUFCMDECUDI(2)",
	OutTemp       => APUFCMDECUDI_OUT(2),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMDECUDI(2),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMDECUDI(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECUDI(3),
	GlitchData    => APUFCMDECUDI3_GlitchData,
	OutSignalName => "APUFCMDECUDI(3)",
	OutTemp       => APUFCMDECUDI_OUT(3),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMDECUDI(3),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMDECUDI(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMDECUDIVALID,
	GlitchData    => APUFCMDECUDIVALID_GlitchData,
	OutSignalName => "APUFCMDECUDIVALID",
	OutTemp       => APUFCMDECUDIVALID_OUT,
	Paths         => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMDECUDIVALID,TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMDECUDIVALID, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMENDIAN,
	GlitchData    => APUFCMENDIAN_GlitchData,
	OutSignalName => "APUFCMENDIAN",
	OutTemp       => APUFCMENDIAN_OUT,
	Paths         => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMENDIAN,TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMENDIAN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMFLUSH,
	GlitchData    => APUFCMFLUSH_GlitchData,
	OutSignalName => "APUFCMFLUSH",
	OutTemp       => APUFCMFLUSH_OUT,
	Paths         => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMFLUSH,TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMFLUSH, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(0),
	GlitchData    => APUFCMINSTRUCTION0_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(0)",
	OutTemp       => APUFCMINSTRUCTION_OUT(0),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(0),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(1),
	GlitchData    => APUFCMINSTRUCTION1_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(1)",
	OutTemp       => APUFCMINSTRUCTION_OUT(1),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(1),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(2),
	GlitchData    => APUFCMINSTRUCTION2_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(2)",
	OutTemp       => APUFCMINSTRUCTION_OUT(2),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(2),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(3),
	GlitchData    => APUFCMINSTRUCTION3_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(3)",
	OutTemp       => APUFCMINSTRUCTION_OUT(3),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(3),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(4),
	GlitchData    => APUFCMINSTRUCTION4_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(4)",
	OutTemp       => APUFCMINSTRUCTION_OUT(4),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(4),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(5),
	GlitchData    => APUFCMINSTRUCTION5_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(5)",
	OutTemp       => APUFCMINSTRUCTION_OUT(5),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(5),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(6),
	GlitchData    => APUFCMINSTRUCTION6_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(6)",
	OutTemp       => APUFCMINSTRUCTION_OUT(6),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(6),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(7),
	GlitchData    => APUFCMINSTRUCTION7_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(7)",
	OutTemp       => APUFCMINSTRUCTION_OUT(7),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(7),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(8),
	GlitchData    => APUFCMINSTRUCTION8_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(8)",
	OutTemp       => APUFCMINSTRUCTION_OUT(8),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(8),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(9),
	GlitchData    => APUFCMINSTRUCTION9_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(9)",
	OutTemp       => APUFCMINSTRUCTION_OUT(9),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(9),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(10),
	GlitchData    => APUFCMINSTRUCTION10_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(10)",
	OutTemp       => APUFCMINSTRUCTION_OUT(10),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(10),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(11),
	GlitchData    => APUFCMINSTRUCTION11_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(11)",
	OutTemp       => APUFCMINSTRUCTION_OUT(11),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(11),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(12),
	GlitchData    => APUFCMINSTRUCTION12_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(12)",
	OutTemp       => APUFCMINSTRUCTION_OUT(12),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(12),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(13),
	GlitchData    => APUFCMINSTRUCTION13_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(13)",
	OutTemp       => APUFCMINSTRUCTION_OUT(13),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(13),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(14),
	GlitchData    => APUFCMINSTRUCTION14_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(14)",
	OutTemp       => APUFCMINSTRUCTION_OUT(14),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(14),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(15),
	GlitchData    => APUFCMINSTRUCTION15_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(15)",
	OutTemp       => APUFCMINSTRUCTION_OUT(15),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(15),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(16),
	GlitchData    => APUFCMINSTRUCTION16_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(16)",
	OutTemp       => APUFCMINSTRUCTION_OUT(16),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(16),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(17),
	GlitchData    => APUFCMINSTRUCTION17_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(17)",
	OutTemp       => APUFCMINSTRUCTION_OUT(17),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(17),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(18),
	GlitchData    => APUFCMINSTRUCTION18_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(18)",
	OutTemp       => APUFCMINSTRUCTION_OUT(18),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(18),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(19),
	GlitchData    => APUFCMINSTRUCTION19_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(19)",
	OutTemp       => APUFCMINSTRUCTION_OUT(19),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(19),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(20),
	GlitchData    => APUFCMINSTRUCTION20_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(20)",
	OutTemp       => APUFCMINSTRUCTION_OUT(20),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(20),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(21),
	GlitchData    => APUFCMINSTRUCTION21_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(21)",
	OutTemp       => APUFCMINSTRUCTION_OUT(21),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(21),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(22),
	GlitchData    => APUFCMINSTRUCTION22_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(22)",
	OutTemp       => APUFCMINSTRUCTION_OUT(22),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(22),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(23),
	GlitchData    => APUFCMINSTRUCTION23_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(23)",
	OutTemp       => APUFCMINSTRUCTION_OUT(23),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(23),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(24),
	GlitchData    => APUFCMINSTRUCTION24_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(24)",
	OutTemp       => APUFCMINSTRUCTION_OUT(24),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(24),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(25),
	GlitchData    => APUFCMINSTRUCTION25_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(25)",
	OutTemp       => APUFCMINSTRUCTION_OUT(25),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(25),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(26),
	GlitchData    => APUFCMINSTRUCTION26_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(26)",
	OutTemp       => APUFCMINSTRUCTION_OUT(26),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(26),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(27),
	GlitchData    => APUFCMINSTRUCTION27_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(27)",
	OutTemp       => APUFCMINSTRUCTION_OUT(27),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(27),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(28),
	GlitchData    => APUFCMINSTRUCTION28_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(28)",
	OutTemp       => APUFCMINSTRUCTION_OUT(28),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(28),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(29),
	GlitchData    => APUFCMINSTRUCTION29_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(29)",
	OutTemp       => APUFCMINSTRUCTION_OUT(29),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(29),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(30),
	GlitchData    => APUFCMINSTRUCTION30_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(30)",
	OutTemp       => APUFCMINSTRUCTION_OUT(30),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(30),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRUCTION(31),
	GlitchData    => APUFCMINSTRUCTION31_GlitchData,
	OutSignalName => "APUFCMINSTRUCTION(31)",
	OutTemp       => APUFCMINSTRUCTION_OUT(31),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRUCTION(31),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRUCTION(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMINSTRVALID,
	GlitchData    => APUFCMINSTRVALID_GlitchData,
	OutSignalName => "APUFCMINSTRVALID",
	OutTemp       => APUFCMINSTRVALID_OUT,
	Paths         => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMINSTRVALID,TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMINSTRVALID, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADBYTEADDR(0),
	GlitchData    => APUFCMLOADBYTEADDR0_GlitchData,
	OutSignalName => "APUFCMLOADBYTEADDR(0)",
	OutTemp       => APUFCMLOADBYTEADDR_OUT(0),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADBYTEADDR(0),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADBYTEADDR(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADBYTEADDR(1),
	GlitchData    => APUFCMLOADBYTEADDR1_GlitchData,
	OutSignalName => "APUFCMLOADBYTEADDR(1)",
	OutTemp       => APUFCMLOADBYTEADDR_OUT(1),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADBYTEADDR(1),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADBYTEADDR(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADBYTEADDR(2),
	GlitchData    => APUFCMLOADBYTEADDR2_GlitchData,
	OutSignalName => "APUFCMLOADBYTEADDR(2)",
	OutTemp       => APUFCMLOADBYTEADDR_OUT(2),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADBYTEADDR(2),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADBYTEADDR(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADBYTEADDR(3),
	GlitchData    => APUFCMLOADBYTEADDR3_GlitchData,
	OutSignalName => "APUFCMLOADBYTEADDR(3)",
	OutTemp       => APUFCMLOADBYTEADDR_OUT(3),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADBYTEADDR(3),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADBYTEADDR(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(0),
	GlitchData    => APUFCMLOADDATA0_GlitchData,
	OutSignalName => "APUFCMLOADDATA(0)",
	OutTemp       => APUFCMLOADDATA_OUT(0),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(0),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(1),
	GlitchData    => APUFCMLOADDATA1_GlitchData,
	OutSignalName => "APUFCMLOADDATA(1)",
	OutTemp       => APUFCMLOADDATA_OUT(1),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(1),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(2),
	GlitchData    => APUFCMLOADDATA2_GlitchData,
	OutSignalName => "APUFCMLOADDATA(2)",
	OutTemp       => APUFCMLOADDATA_OUT(2),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(2),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(3),
	GlitchData    => APUFCMLOADDATA3_GlitchData,
	OutSignalName => "APUFCMLOADDATA(3)",
	OutTemp       => APUFCMLOADDATA_OUT(3),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(3),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(4),
	GlitchData    => APUFCMLOADDATA4_GlitchData,
	OutSignalName => "APUFCMLOADDATA(4)",
	OutTemp       => APUFCMLOADDATA_OUT(4),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(4),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(5),
	GlitchData    => APUFCMLOADDATA5_GlitchData,
	OutSignalName => "APUFCMLOADDATA(5)",
	OutTemp       => APUFCMLOADDATA_OUT(5),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(5),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(6),
	GlitchData    => APUFCMLOADDATA6_GlitchData,
	OutSignalName => "APUFCMLOADDATA(6)",
	OutTemp       => APUFCMLOADDATA_OUT(6),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(6),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(7),
	GlitchData    => APUFCMLOADDATA7_GlitchData,
	OutSignalName => "APUFCMLOADDATA(7)",
	OutTemp       => APUFCMLOADDATA_OUT(7),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(7),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(8),
	GlitchData    => APUFCMLOADDATA8_GlitchData,
	OutSignalName => "APUFCMLOADDATA(8)",
	OutTemp       => APUFCMLOADDATA_OUT(8),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(8),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(9),
	GlitchData    => APUFCMLOADDATA9_GlitchData,
	OutSignalName => "APUFCMLOADDATA(9)",
	OutTemp       => APUFCMLOADDATA_OUT(9),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(9),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(10),
	GlitchData    => APUFCMLOADDATA10_GlitchData,
	OutSignalName => "APUFCMLOADDATA(10)",
	OutTemp       => APUFCMLOADDATA_OUT(10),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(10),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(11),
	GlitchData    => APUFCMLOADDATA11_GlitchData,
	OutSignalName => "APUFCMLOADDATA(11)",
	OutTemp       => APUFCMLOADDATA_OUT(11),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(11),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(12),
	GlitchData    => APUFCMLOADDATA12_GlitchData,
	OutSignalName => "APUFCMLOADDATA(12)",
	OutTemp       => APUFCMLOADDATA_OUT(12),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(12),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(13),
	GlitchData    => APUFCMLOADDATA13_GlitchData,
	OutSignalName => "APUFCMLOADDATA(13)",
	OutTemp       => APUFCMLOADDATA_OUT(13),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(13),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(14),
	GlitchData    => APUFCMLOADDATA14_GlitchData,
	OutSignalName => "APUFCMLOADDATA(14)",
	OutTemp       => APUFCMLOADDATA_OUT(14),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(14),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(15),
	GlitchData    => APUFCMLOADDATA15_GlitchData,
	OutSignalName => "APUFCMLOADDATA(15)",
	OutTemp       => APUFCMLOADDATA_OUT(15),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(15),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(16),
	GlitchData    => APUFCMLOADDATA16_GlitchData,
	OutSignalName => "APUFCMLOADDATA(16)",
	OutTemp       => APUFCMLOADDATA_OUT(16),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(16),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(17),
	GlitchData    => APUFCMLOADDATA17_GlitchData,
	OutSignalName => "APUFCMLOADDATA(17)",
	OutTemp       => APUFCMLOADDATA_OUT(17),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(17),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(18),
	GlitchData    => APUFCMLOADDATA18_GlitchData,
	OutSignalName => "APUFCMLOADDATA(18)",
	OutTemp       => APUFCMLOADDATA_OUT(18),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(18),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(19),
	GlitchData    => APUFCMLOADDATA19_GlitchData,
	OutSignalName => "APUFCMLOADDATA(19)",
	OutTemp       => APUFCMLOADDATA_OUT(19),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(19),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(20),
	GlitchData    => APUFCMLOADDATA20_GlitchData,
	OutSignalName => "APUFCMLOADDATA(20)",
	OutTemp       => APUFCMLOADDATA_OUT(20),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(20),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(21),
	GlitchData    => APUFCMLOADDATA21_GlitchData,
	OutSignalName => "APUFCMLOADDATA(21)",
	OutTemp       => APUFCMLOADDATA_OUT(21),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(21),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(22),
	GlitchData    => APUFCMLOADDATA22_GlitchData,
	OutSignalName => "APUFCMLOADDATA(22)",
	OutTemp       => APUFCMLOADDATA_OUT(22),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(22),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(23),
	GlitchData    => APUFCMLOADDATA23_GlitchData,
	OutSignalName => "APUFCMLOADDATA(23)",
	OutTemp       => APUFCMLOADDATA_OUT(23),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(23),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(24),
	GlitchData    => APUFCMLOADDATA24_GlitchData,
	OutSignalName => "APUFCMLOADDATA(24)",
	OutTemp       => APUFCMLOADDATA_OUT(24),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(24),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(25),
	GlitchData    => APUFCMLOADDATA25_GlitchData,
	OutSignalName => "APUFCMLOADDATA(25)",
	OutTemp       => APUFCMLOADDATA_OUT(25),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(25),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(26),
	GlitchData    => APUFCMLOADDATA26_GlitchData,
	OutSignalName => "APUFCMLOADDATA(26)",
	OutTemp       => APUFCMLOADDATA_OUT(26),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(26),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(27),
	GlitchData    => APUFCMLOADDATA27_GlitchData,
	OutSignalName => "APUFCMLOADDATA(27)",
	OutTemp       => APUFCMLOADDATA_OUT(27),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(27),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(28),
	GlitchData    => APUFCMLOADDATA28_GlitchData,
	OutSignalName => "APUFCMLOADDATA(28)",
	OutTemp       => APUFCMLOADDATA_OUT(28),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(28),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(29),
	GlitchData    => APUFCMLOADDATA29_GlitchData,
	OutSignalName => "APUFCMLOADDATA(29)",
	OutTemp       => APUFCMLOADDATA_OUT(29),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(29),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(30),
	GlitchData    => APUFCMLOADDATA30_GlitchData,
	OutSignalName => "APUFCMLOADDATA(30)",
	OutTemp       => APUFCMLOADDATA_OUT(30),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(30),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(31),
	GlitchData    => APUFCMLOADDATA31_GlitchData,
	OutSignalName => "APUFCMLOADDATA(31)",
	OutTemp       => APUFCMLOADDATA_OUT(31),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(31),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(32),
	GlitchData    => APUFCMLOADDATA32_GlitchData,
	OutSignalName => "APUFCMLOADDATA(32)",
	OutTemp       => APUFCMLOADDATA_OUT(32),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(32),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(32), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(33),
	GlitchData    => APUFCMLOADDATA33_GlitchData,
	OutSignalName => "APUFCMLOADDATA(33)",
	OutTemp       => APUFCMLOADDATA_OUT(33),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(33),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(33), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(34),
	GlitchData    => APUFCMLOADDATA34_GlitchData,
	OutSignalName => "APUFCMLOADDATA(34)",
	OutTemp       => APUFCMLOADDATA_OUT(34),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(34),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(34), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(35),
	GlitchData    => APUFCMLOADDATA35_GlitchData,
	OutSignalName => "APUFCMLOADDATA(35)",
	OutTemp       => APUFCMLOADDATA_OUT(35),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(35),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(35), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(36),
	GlitchData    => APUFCMLOADDATA36_GlitchData,
	OutSignalName => "APUFCMLOADDATA(36)",
	OutTemp       => APUFCMLOADDATA_OUT(36),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(36),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(36), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(37),
	GlitchData    => APUFCMLOADDATA37_GlitchData,
	OutSignalName => "APUFCMLOADDATA(37)",
	OutTemp       => APUFCMLOADDATA_OUT(37),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(37),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(37), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(38),
	GlitchData    => APUFCMLOADDATA38_GlitchData,
	OutSignalName => "APUFCMLOADDATA(38)",
	OutTemp       => APUFCMLOADDATA_OUT(38),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(38),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(38), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(39),
	GlitchData    => APUFCMLOADDATA39_GlitchData,
	OutSignalName => "APUFCMLOADDATA(39)",
	OutTemp       => APUFCMLOADDATA_OUT(39),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(39),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(39), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(40),
	GlitchData    => APUFCMLOADDATA40_GlitchData,
	OutSignalName => "APUFCMLOADDATA(40)",
	OutTemp       => APUFCMLOADDATA_OUT(40),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(40),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(40), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(41),
	GlitchData    => APUFCMLOADDATA41_GlitchData,
	OutSignalName => "APUFCMLOADDATA(41)",
	OutTemp       => APUFCMLOADDATA_OUT(41),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(41),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(41), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(42),
	GlitchData    => APUFCMLOADDATA42_GlitchData,
	OutSignalName => "APUFCMLOADDATA(42)",
	OutTemp       => APUFCMLOADDATA_OUT(42),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(42),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(42), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(43),
	GlitchData    => APUFCMLOADDATA43_GlitchData,
	OutSignalName => "APUFCMLOADDATA(43)",
	OutTemp       => APUFCMLOADDATA_OUT(43),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(43),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(43), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(44),
	GlitchData    => APUFCMLOADDATA44_GlitchData,
	OutSignalName => "APUFCMLOADDATA(44)",
	OutTemp       => APUFCMLOADDATA_OUT(44),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(44),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(44), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(45),
	GlitchData    => APUFCMLOADDATA45_GlitchData,
	OutSignalName => "APUFCMLOADDATA(45)",
	OutTemp       => APUFCMLOADDATA_OUT(45),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(45),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(45), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(46),
	GlitchData    => APUFCMLOADDATA46_GlitchData,
	OutSignalName => "APUFCMLOADDATA(46)",
	OutTemp       => APUFCMLOADDATA_OUT(46),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(46),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(46), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(47),
	GlitchData    => APUFCMLOADDATA47_GlitchData,
	OutSignalName => "APUFCMLOADDATA(47)",
	OutTemp       => APUFCMLOADDATA_OUT(47),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(47),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(47), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(48),
	GlitchData    => APUFCMLOADDATA48_GlitchData,
	OutSignalName => "APUFCMLOADDATA(48)",
	OutTemp       => APUFCMLOADDATA_OUT(48),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(48),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(48), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(49),
	GlitchData    => APUFCMLOADDATA49_GlitchData,
	OutSignalName => "APUFCMLOADDATA(49)",
	OutTemp       => APUFCMLOADDATA_OUT(49),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(49),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(49), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(50),
	GlitchData    => APUFCMLOADDATA50_GlitchData,
	OutSignalName => "APUFCMLOADDATA(50)",
	OutTemp       => APUFCMLOADDATA_OUT(50),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(50),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(50), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(51),
	GlitchData    => APUFCMLOADDATA51_GlitchData,
	OutSignalName => "APUFCMLOADDATA(51)",
	OutTemp       => APUFCMLOADDATA_OUT(51),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(51),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(51), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(52),
	GlitchData    => APUFCMLOADDATA52_GlitchData,
	OutSignalName => "APUFCMLOADDATA(52)",
	OutTemp       => APUFCMLOADDATA_OUT(52),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(52),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(52), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(53),
	GlitchData    => APUFCMLOADDATA53_GlitchData,
	OutSignalName => "APUFCMLOADDATA(53)",
	OutTemp       => APUFCMLOADDATA_OUT(53),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(53),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(53), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(54),
	GlitchData    => APUFCMLOADDATA54_GlitchData,
	OutSignalName => "APUFCMLOADDATA(54)",
	OutTemp       => APUFCMLOADDATA_OUT(54),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(54),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(54), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(55),
	GlitchData    => APUFCMLOADDATA55_GlitchData,
	OutSignalName => "APUFCMLOADDATA(55)",
	OutTemp       => APUFCMLOADDATA_OUT(55),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(55),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(55), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(56),
	GlitchData    => APUFCMLOADDATA56_GlitchData,
	OutSignalName => "APUFCMLOADDATA(56)",
	OutTemp       => APUFCMLOADDATA_OUT(56),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(56),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(56), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(57),
	GlitchData    => APUFCMLOADDATA57_GlitchData,
	OutSignalName => "APUFCMLOADDATA(57)",
	OutTemp       => APUFCMLOADDATA_OUT(57),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(57),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(57), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(58),
	GlitchData    => APUFCMLOADDATA58_GlitchData,
	OutSignalName => "APUFCMLOADDATA(58)",
	OutTemp       => APUFCMLOADDATA_OUT(58),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(58),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(58), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(59),
	GlitchData    => APUFCMLOADDATA59_GlitchData,
	OutSignalName => "APUFCMLOADDATA(59)",
	OutTemp       => APUFCMLOADDATA_OUT(59),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(59),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(59), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(60),
	GlitchData    => APUFCMLOADDATA60_GlitchData,
	OutSignalName => "APUFCMLOADDATA(60)",
	OutTemp       => APUFCMLOADDATA_OUT(60),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(60),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(60), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(61),
	GlitchData    => APUFCMLOADDATA61_GlitchData,
	OutSignalName => "APUFCMLOADDATA(61)",
	OutTemp       => APUFCMLOADDATA_OUT(61),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(61),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(61), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(62),
	GlitchData    => APUFCMLOADDATA62_GlitchData,
	OutSignalName => "APUFCMLOADDATA(62)",
	OutTemp       => APUFCMLOADDATA_OUT(62),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(62),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(62), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(63),
	GlitchData    => APUFCMLOADDATA63_GlitchData,
	OutSignalName => "APUFCMLOADDATA(63)",
	OutTemp       => APUFCMLOADDATA_OUT(63),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(63),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(63), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(64),
	GlitchData    => APUFCMLOADDATA64_GlitchData,
	OutSignalName => "APUFCMLOADDATA(64)",
	OutTemp       => APUFCMLOADDATA_OUT(64),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(64),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(64), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(65),
	GlitchData    => APUFCMLOADDATA65_GlitchData,
	OutSignalName => "APUFCMLOADDATA(65)",
	OutTemp       => APUFCMLOADDATA_OUT(65),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(65),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(65), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(66),
	GlitchData    => APUFCMLOADDATA66_GlitchData,
	OutSignalName => "APUFCMLOADDATA(66)",
	OutTemp       => APUFCMLOADDATA_OUT(66),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(66),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(66), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(67),
	GlitchData    => APUFCMLOADDATA67_GlitchData,
	OutSignalName => "APUFCMLOADDATA(67)",
	OutTemp       => APUFCMLOADDATA_OUT(67),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(67),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(67), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(68),
	GlitchData    => APUFCMLOADDATA68_GlitchData,
	OutSignalName => "APUFCMLOADDATA(68)",
	OutTemp       => APUFCMLOADDATA_OUT(68),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(68),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(68), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(69),
	GlitchData    => APUFCMLOADDATA69_GlitchData,
	OutSignalName => "APUFCMLOADDATA(69)",
	OutTemp       => APUFCMLOADDATA_OUT(69),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(69),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(69), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(70),
	GlitchData    => APUFCMLOADDATA70_GlitchData,
	OutSignalName => "APUFCMLOADDATA(70)",
	OutTemp       => APUFCMLOADDATA_OUT(70),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(70),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(70), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(71),
	GlitchData    => APUFCMLOADDATA71_GlitchData,
	OutSignalName => "APUFCMLOADDATA(71)",
	OutTemp       => APUFCMLOADDATA_OUT(71),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(71),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(71), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(72),
	GlitchData    => APUFCMLOADDATA72_GlitchData,
	OutSignalName => "APUFCMLOADDATA(72)",
	OutTemp       => APUFCMLOADDATA_OUT(72),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(72),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(72), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(73),
	GlitchData    => APUFCMLOADDATA73_GlitchData,
	OutSignalName => "APUFCMLOADDATA(73)",
	OutTemp       => APUFCMLOADDATA_OUT(73),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(73),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(73), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(74),
	GlitchData    => APUFCMLOADDATA74_GlitchData,
	OutSignalName => "APUFCMLOADDATA(74)",
	OutTemp       => APUFCMLOADDATA_OUT(74),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(74),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(74), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(75),
	GlitchData    => APUFCMLOADDATA75_GlitchData,
	OutSignalName => "APUFCMLOADDATA(75)",
	OutTemp       => APUFCMLOADDATA_OUT(75),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(75),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(75), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(76),
	GlitchData    => APUFCMLOADDATA76_GlitchData,
	OutSignalName => "APUFCMLOADDATA(76)",
	OutTemp       => APUFCMLOADDATA_OUT(76),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(76),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(76), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(77),
	GlitchData    => APUFCMLOADDATA77_GlitchData,
	OutSignalName => "APUFCMLOADDATA(77)",
	OutTemp       => APUFCMLOADDATA_OUT(77),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(77),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(77), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(78),
	GlitchData    => APUFCMLOADDATA78_GlitchData,
	OutSignalName => "APUFCMLOADDATA(78)",
	OutTemp       => APUFCMLOADDATA_OUT(78),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(78),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(78), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(79),
	GlitchData    => APUFCMLOADDATA79_GlitchData,
	OutSignalName => "APUFCMLOADDATA(79)",
	OutTemp       => APUFCMLOADDATA_OUT(79),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(79),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(79), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(80),
	GlitchData    => APUFCMLOADDATA80_GlitchData,
	OutSignalName => "APUFCMLOADDATA(80)",
	OutTemp       => APUFCMLOADDATA_OUT(80),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(80),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(80), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(81),
	GlitchData    => APUFCMLOADDATA81_GlitchData,
	OutSignalName => "APUFCMLOADDATA(81)",
	OutTemp       => APUFCMLOADDATA_OUT(81),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(81),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(81), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(82),
	GlitchData    => APUFCMLOADDATA82_GlitchData,
	OutSignalName => "APUFCMLOADDATA(82)",
	OutTemp       => APUFCMLOADDATA_OUT(82),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(82),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(82), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(83),
	GlitchData    => APUFCMLOADDATA83_GlitchData,
	OutSignalName => "APUFCMLOADDATA(83)",
	OutTemp       => APUFCMLOADDATA_OUT(83),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(83),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(83), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(84),
	GlitchData    => APUFCMLOADDATA84_GlitchData,
	OutSignalName => "APUFCMLOADDATA(84)",
	OutTemp       => APUFCMLOADDATA_OUT(84),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(84),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(84), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(85),
	GlitchData    => APUFCMLOADDATA85_GlitchData,
	OutSignalName => "APUFCMLOADDATA(85)",
	OutTemp       => APUFCMLOADDATA_OUT(85),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(85),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(85), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(86),
	GlitchData    => APUFCMLOADDATA86_GlitchData,
	OutSignalName => "APUFCMLOADDATA(86)",
	OutTemp       => APUFCMLOADDATA_OUT(86),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(86),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(86), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(87),
	GlitchData    => APUFCMLOADDATA87_GlitchData,
	OutSignalName => "APUFCMLOADDATA(87)",
	OutTemp       => APUFCMLOADDATA_OUT(87),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(87),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(87), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(88),
	GlitchData    => APUFCMLOADDATA88_GlitchData,
	OutSignalName => "APUFCMLOADDATA(88)",
	OutTemp       => APUFCMLOADDATA_OUT(88),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(88),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(88), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(89),
	GlitchData    => APUFCMLOADDATA89_GlitchData,
	OutSignalName => "APUFCMLOADDATA(89)",
	OutTemp       => APUFCMLOADDATA_OUT(89),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(89),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(89), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(90),
	GlitchData    => APUFCMLOADDATA90_GlitchData,
	OutSignalName => "APUFCMLOADDATA(90)",
	OutTemp       => APUFCMLOADDATA_OUT(90),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(90),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(90), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(91),
	GlitchData    => APUFCMLOADDATA91_GlitchData,
	OutSignalName => "APUFCMLOADDATA(91)",
	OutTemp       => APUFCMLOADDATA_OUT(91),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(91),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(91), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(92),
	GlitchData    => APUFCMLOADDATA92_GlitchData,
	OutSignalName => "APUFCMLOADDATA(92)",
	OutTemp       => APUFCMLOADDATA_OUT(92),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(92),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(92), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(93),
	GlitchData    => APUFCMLOADDATA93_GlitchData,
	OutSignalName => "APUFCMLOADDATA(93)",
	OutTemp       => APUFCMLOADDATA_OUT(93),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(93),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(93), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(94),
	GlitchData    => APUFCMLOADDATA94_GlitchData,
	OutSignalName => "APUFCMLOADDATA(94)",
	OutTemp       => APUFCMLOADDATA_OUT(94),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(94),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(94), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(95),
	GlitchData    => APUFCMLOADDATA95_GlitchData,
	OutSignalName => "APUFCMLOADDATA(95)",
	OutTemp       => APUFCMLOADDATA_OUT(95),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(95),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(95), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(96),
	GlitchData    => APUFCMLOADDATA96_GlitchData,
	OutSignalName => "APUFCMLOADDATA(96)",
	OutTemp       => APUFCMLOADDATA_OUT(96),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(96),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(96), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(97),
	GlitchData    => APUFCMLOADDATA97_GlitchData,
	OutSignalName => "APUFCMLOADDATA(97)",
	OutTemp       => APUFCMLOADDATA_OUT(97),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(97),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(97), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(98),
	GlitchData    => APUFCMLOADDATA98_GlitchData,
	OutSignalName => "APUFCMLOADDATA(98)",
	OutTemp       => APUFCMLOADDATA_OUT(98),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(98),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(98), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(99),
	GlitchData    => APUFCMLOADDATA99_GlitchData,
	OutSignalName => "APUFCMLOADDATA(99)",
	OutTemp       => APUFCMLOADDATA_OUT(99),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(99),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(99), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(100),
	GlitchData    => APUFCMLOADDATA100_GlitchData,
	OutSignalName => "APUFCMLOADDATA(100)",
	OutTemp       => APUFCMLOADDATA_OUT(100),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(100),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(100), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(101),
	GlitchData    => APUFCMLOADDATA101_GlitchData,
	OutSignalName => "APUFCMLOADDATA(101)",
	OutTemp       => APUFCMLOADDATA_OUT(101),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(101),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(101), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(102),
	GlitchData    => APUFCMLOADDATA102_GlitchData,
	OutSignalName => "APUFCMLOADDATA(102)",
	OutTemp       => APUFCMLOADDATA_OUT(102),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(102),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(102), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(103),
	GlitchData    => APUFCMLOADDATA103_GlitchData,
	OutSignalName => "APUFCMLOADDATA(103)",
	OutTemp       => APUFCMLOADDATA_OUT(103),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(103),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(103), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(104),
	GlitchData    => APUFCMLOADDATA104_GlitchData,
	OutSignalName => "APUFCMLOADDATA(104)",
	OutTemp       => APUFCMLOADDATA_OUT(104),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(104),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(104), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(105),
	GlitchData    => APUFCMLOADDATA105_GlitchData,
	OutSignalName => "APUFCMLOADDATA(105)",
	OutTemp       => APUFCMLOADDATA_OUT(105),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(105),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(105), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(106),
	GlitchData    => APUFCMLOADDATA106_GlitchData,
	OutSignalName => "APUFCMLOADDATA(106)",
	OutTemp       => APUFCMLOADDATA_OUT(106),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(106),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(106), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(107),
	GlitchData    => APUFCMLOADDATA107_GlitchData,
	OutSignalName => "APUFCMLOADDATA(107)",
	OutTemp       => APUFCMLOADDATA_OUT(107),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(107),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(107), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(108),
	GlitchData    => APUFCMLOADDATA108_GlitchData,
	OutSignalName => "APUFCMLOADDATA(108)",
	OutTemp       => APUFCMLOADDATA_OUT(108),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(108),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(108), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(109),
	GlitchData    => APUFCMLOADDATA109_GlitchData,
	OutSignalName => "APUFCMLOADDATA(109)",
	OutTemp       => APUFCMLOADDATA_OUT(109),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(109),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(109), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(110),
	GlitchData    => APUFCMLOADDATA110_GlitchData,
	OutSignalName => "APUFCMLOADDATA(110)",
	OutTemp       => APUFCMLOADDATA_OUT(110),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(110),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(110), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(111),
	GlitchData    => APUFCMLOADDATA111_GlitchData,
	OutSignalName => "APUFCMLOADDATA(111)",
	OutTemp       => APUFCMLOADDATA_OUT(111),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(111),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(111), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(112),
	GlitchData    => APUFCMLOADDATA112_GlitchData,
	OutSignalName => "APUFCMLOADDATA(112)",
	OutTemp       => APUFCMLOADDATA_OUT(112),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(112),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(112), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(113),
	GlitchData    => APUFCMLOADDATA113_GlitchData,
	OutSignalName => "APUFCMLOADDATA(113)",
	OutTemp       => APUFCMLOADDATA_OUT(113),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(113),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(113), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(114),
	GlitchData    => APUFCMLOADDATA114_GlitchData,
	OutSignalName => "APUFCMLOADDATA(114)",
	OutTemp       => APUFCMLOADDATA_OUT(114),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(114),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(114), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(115),
	GlitchData    => APUFCMLOADDATA115_GlitchData,
	OutSignalName => "APUFCMLOADDATA(115)",
	OutTemp       => APUFCMLOADDATA_OUT(115),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(115),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(115), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(116),
	GlitchData    => APUFCMLOADDATA116_GlitchData,
	OutSignalName => "APUFCMLOADDATA(116)",
	OutTemp       => APUFCMLOADDATA_OUT(116),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(116),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(116), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(117),
	GlitchData    => APUFCMLOADDATA117_GlitchData,
	OutSignalName => "APUFCMLOADDATA(117)",
	OutTemp       => APUFCMLOADDATA_OUT(117),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(117),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(117), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(118),
	GlitchData    => APUFCMLOADDATA118_GlitchData,
	OutSignalName => "APUFCMLOADDATA(118)",
	OutTemp       => APUFCMLOADDATA_OUT(118),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(118),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(118), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(119),
	GlitchData    => APUFCMLOADDATA119_GlitchData,
	OutSignalName => "APUFCMLOADDATA(119)",
	OutTemp       => APUFCMLOADDATA_OUT(119),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(119),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(119), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(120),
	GlitchData    => APUFCMLOADDATA120_GlitchData,
	OutSignalName => "APUFCMLOADDATA(120)",
	OutTemp       => APUFCMLOADDATA_OUT(120),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(120),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(120), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(121),
	GlitchData    => APUFCMLOADDATA121_GlitchData,
	OutSignalName => "APUFCMLOADDATA(121)",
	OutTemp       => APUFCMLOADDATA_OUT(121),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(121),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(121), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(122),
	GlitchData    => APUFCMLOADDATA122_GlitchData,
	OutSignalName => "APUFCMLOADDATA(122)",
	OutTemp       => APUFCMLOADDATA_OUT(122),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(122),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(122), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(123),
	GlitchData    => APUFCMLOADDATA123_GlitchData,
	OutSignalName => "APUFCMLOADDATA(123)",
	OutTemp       => APUFCMLOADDATA_OUT(123),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(123),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(123), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(124),
	GlitchData    => APUFCMLOADDATA124_GlitchData,
	OutSignalName => "APUFCMLOADDATA(124)",
	OutTemp       => APUFCMLOADDATA_OUT(124),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(124),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(124), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(125),
	GlitchData    => APUFCMLOADDATA125_GlitchData,
	OutSignalName => "APUFCMLOADDATA(125)",
	OutTemp       => APUFCMLOADDATA_OUT(125),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(125),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(125), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(126),
	GlitchData    => APUFCMLOADDATA126_GlitchData,
	OutSignalName => "APUFCMLOADDATA(126)",
	OutTemp       => APUFCMLOADDATA_OUT(126),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(126),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(126), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDATA(127),
	GlitchData    => APUFCMLOADDATA127_GlitchData,
	OutSignalName => "APUFCMLOADDATA(127)",
	OutTemp       => APUFCMLOADDATA_OUT(127),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDATA(127),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDATA(127), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMLOADDVALID,
	GlitchData    => APUFCMLOADDVALID_GlitchData,
	OutSignalName => "APUFCMLOADDVALID",
	OutTemp       => APUFCMLOADDVALID_OUT,
	Paths         => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMLOADDVALID,TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMLOADDVALID, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMMSRFE0,
	GlitchData    => APUFCMMSRFE0_GlitchData,
	OutSignalName => "APUFCMMSRFE0",
	OutTemp       => APUFCMMSRFE0_OUT,
	Paths         => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMMSRFE0,TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMMSRFE0, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMMSRFE1,
	GlitchData    => APUFCMMSRFE1_GlitchData,
	OutSignalName => "APUFCMMSRFE1",
	OutTemp       => APUFCMMSRFE1_OUT,
	Paths         => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMMSRFE1,TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMMSRFE1, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMNEXTINSTRREADY,
	GlitchData    => APUFCMNEXTINSTRREADY_GlitchData,
	OutSignalName => "APUFCMNEXTINSTRREADY",
	OutTemp       => APUFCMNEXTINSTRREADY_OUT,
	Paths         => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMNEXTINSTRREADY,TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMNEXTINSTRREADY, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMOPERANDVALID,
	GlitchData    => APUFCMOPERANDVALID_GlitchData,
	OutSignalName => "APUFCMOPERANDVALID",
	OutTemp       => APUFCMOPERANDVALID_OUT,
	Paths         => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMOPERANDVALID,TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMOPERANDVALID, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(0),
	GlitchData    => APUFCMRADATA0_GlitchData,
	OutSignalName => "APUFCMRADATA(0)",
	OutTemp       => APUFCMRADATA_OUT(0),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(0),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(1),
	GlitchData    => APUFCMRADATA1_GlitchData,
	OutSignalName => "APUFCMRADATA(1)",
	OutTemp       => APUFCMRADATA_OUT(1),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(1),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(2),
	GlitchData    => APUFCMRADATA2_GlitchData,
	OutSignalName => "APUFCMRADATA(2)",
	OutTemp       => APUFCMRADATA_OUT(2),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(2),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(3),
	GlitchData    => APUFCMRADATA3_GlitchData,
	OutSignalName => "APUFCMRADATA(3)",
	OutTemp       => APUFCMRADATA_OUT(3),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(3),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(4),
	GlitchData    => APUFCMRADATA4_GlitchData,
	OutSignalName => "APUFCMRADATA(4)",
	OutTemp       => APUFCMRADATA_OUT(4),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(4),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(5),
	GlitchData    => APUFCMRADATA5_GlitchData,
	OutSignalName => "APUFCMRADATA(5)",
	OutTemp       => APUFCMRADATA_OUT(5),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(5),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(6),
	GlitchData    => APUFCMRADATA6_GlitchData,
	OutSignalName => "APUFCMRADATA(6)",
	OutTemp       => APUFCMRADATA_OUT(6),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(6),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(7),
	GlitchData    => APUFCMRADATA7_GlitchData,
	OutSignalName => "APUFCMRADATA(7)",
	OutTemp       => APUFCMRADATA_OUT(7),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(7),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(8),
	GlitchData    => APUFCMRADATA8_GlitchData,
	OutSignalName => "APUFCMRADATA(8)",
	OutTemp       => APUFCMRADATA_OUT(8),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(8),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(9),
	GlitchData    => APUFCMRADATA9_GlitchData,
	OutSignalName => "APUFCMRADATA(9)",
	OutTemp       => APUFCMRADATA_OUT(9),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(9),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(10),
	GlitchData    => APUFCMRADATA10_GlitchData,
	OutSignalName => "APUFCMRADATA(10)",
	OutTemp       => APUFCMRADATA_OUT(10),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(10),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(11),
	GlitchData    => APUFCMRADATA11_GlitchData,
	OutSignalName => "APUFCMRADATA(11)",
	OutTemp       => APUFCMRADATA_OUT(11),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(11),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(12),
	GlitchData    => APUFCMRADATA12_GlitchData,
	OutSignalName => "APUFCMRADATA(12)",
	OutTemp       => APUFCMRADATA_OUT(12),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(12),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(13),
	GlitchData    => APUFCMRADATA13_GlitchData,
	OutSignalName => "APUFCMRADATA(13)",
	OutTemp       => APUFCMRADATA_OUT(13),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(13),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(14),
	GlitchData    => APUFCMRADATA14_GlitchData,
	OutSignalName => "APUFCMRADATA(14)",
	OutTemp       => APUFCMRADATA_OUT(14),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(14),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(15),
	GlitchData    => APUFCMRADATA15_GlitchData,
	OutSignalName => "APUFCMRADATA(15)",
	OutTemp       => APUFCMRADATA_OUT(15),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(15),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(16),
	GlitchData    => APUFCMRADATA16_GlitchData,
	OutSignalName => "APUFCMRADATA(16)",
	OutTemp       => APUFCMRADATA_OUT(16),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(16),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(17),
	GlitchData    => APUFCMRADATA17_GlitchData,
	OutSignalName => "APUFCMRADATA(17)",
	OutTemp       => APUFCMRADATA_OUT(17),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(17),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(18),
	GlitchData    => APUFCMRADATA18_GlitchData,
	OutSignalName => "APUFCMRADATA(18)",
	OutTemp       => APUFCMRADATA_OUT(18),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(18),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(19),
	GlitchData    => APUFCMRADATA19_GlitchData,
	OutSignalName => "APUFCMRADATA(19)",
	OutTemp       => APUFCMRADATA_OUT(19),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(19),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(20),
	GlitchData    => APUFCMRADATA20_GlitchData,
	OutSignalName => "APUFCMRADATA(20)",
	OutTemp       => APUFCMRADATA_OUT(20),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(20),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(21),
	GlitchData    => APUFCMRADATA21_GlitchData,
	OutSignalName => "APUFCMRADATA(21)",
	OutTemp       => APUFCMRADATA_OUT(21),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(21),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(22),
	GlitchData    => APUFCMRADATA22_GlitchData,
	OutSignalName => "APUFCMRADATA(22)",
	OutTemp       => APUFCMRADATA_OUT(22),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(22),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(23),
	GlitchData    => APUFCMRADATA23_GlitchData,
	OutSignalName => "APUFCMRADATA(23)",
	OutTemp       => APUFCMRADATA_OUT(23),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(23),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(24),
	GlitchData    => APUFCMRADATA24_GlitchData,
	OutSignalName => "APUFCMRADATA(24)",
	OutTemp       => APUFCMRADATA_OUT(24),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(24),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(25),
	GlitchData    => APUFCMRADATA25_GlitchData,
	OutSignalName => "APUFCMRADATA(25)",
	OutTemp       => APUFCMRADATA_OUT(25),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(25),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(26),
	GlitchData    => APUFCMRADATA26_GlitchData,
	OutSignalName => "APUFCMRADATA(26)",
	OutTemp       => APUFCMRADATA_OUT(26),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(26),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(27),
	GlitchData    => APUFCMRADATA27_GlitchData,
	OutSignalName => "APUFCMRADATA(27)",
	OutTemp       => APUFCMRADATA_OUT(27),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(27),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(28),
	GlitchData    => APUFCMRADATA28_GlitchData,
	OutSignalName => "APUFCMRADATA(28)",
	OutTemp       => APUFCMRADATA_OUT(28),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(28),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(29),
	GlitchData    => APUFCMRADATA29_GlitchData,
	OutSignalName => "APUFCMRADATA(29)",
	OutTemp       => APUFCMRADATA_OUT(29),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(29),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(30),
	GlitchData    => APUFCMRADATA30_GlitchData,
	OutSignalName => "APUFCMRADATA(30)",
	OutTemp       => APUFCMRADATA_OUT(30),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(30),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRADATA(31),
	GlitchData    => APUFCMRADATA31_GlitchData,
	OutSignalName => "APUFCMRADATA(31)",
	OutTemp       => APUFCMRADATA_OUT(31),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRADATA(31),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRADATA(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(0),
	GlitchData    => APUFCMRBDATA0_GlitchData,
	OutSignalName => "APUFCMRBDATA(0)",
	OutTemp       => APUFCMRBDATA_OUT(0),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(0),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(1),
	GlitchData    => APUFCMRBDATA1_GlitchData,
	OutSignalName => "APUFCMRBDATA(1)",
	OutTemp       => APUFCMRBDATA_OUT(1),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(1),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(2),
	GlitchData    => APUFCMRBDATA2_GlitchData,
	OutSignalName => "APUFCMRBDATA(2)",
	OutTemp       => APUFCMRBDATA_OUT(2),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(2),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(3),
	GlitchData    => APUFCMRBDATA3_GlitchData,
	OutSignalName => "APUFCMRBDATA(3)",
	OutTemp       => APUFCMRBDATA_OUT(3),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(3),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(4),
	GlitchData    => APUFCMRBDATA4_GlitchData,
	OutSignalName => "APUFCMRBDATA(4)",
	OutTemp       => APUFCMRBDATA_OUT(4),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(4),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(5),
	GlitchData    => APUFCMRBDATA5_GlitchData,
	OutSignalName => "APUFCMRBDATA(5)",
	OutTemp       => APUFCMRBDATA_OUT(5),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(5),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(6),
	GlitchData    => APUFCMRBDATA6_GlitchData,
	OutSignalName => "APUFCMRBDATA(6)",
	OutTemp       => APUFCMRBDATA_OUT(6),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(6),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(7),
	GlitchData    => APUFCMRBDATA7_GlitchData,
	OutSignalName => "APUFCMRBDATA(7)",
	OutTemp       => APUFCMRBDATA_OUT(7),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(7),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(8),
	GlitchData    => APUFCMRBDATA8_GlitchData,
	OutSignalName => "APUFCMRBDATA(8)",
	OutTemp       => APUFCMRBDATA_OUT(8),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(8),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(9),
	GlitchData    => APUFCMRBDATA9_GlitchData,
	OutSignalName => "APUFCMRBDATA(9)",
	OutTemp       => APUFCMRBDATA_OUT(9),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(9),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(10),
	GlitchData    => APUFCMRBDATA10_GlitchData,
	OutSignalName => "APUFCMRBDATA(10)",
	OutTemp       => APUFCMRBDATA_OUT(10),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(10),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(11),
	GlitchData    => APUFCMRBDATA11_GlitchData,
	OutSignalName => "APUFCMRBDATA(11)",
	OutTemp       => APUFCMRBDATA_OUT(11),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(11),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(12),
	GlitchData    => APUFCMRBDATA12_GlitchData,
	OutSignalName => "APUFCMRBDATA(12)",
	OutTemp       => APUFCMRBDATA_OUT(12),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(12),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(13),
	GlitchData    => APUFCMRBDATA13_GlitchData,
	OutSignalName => "APUFCMRBDATA(13)",
	OutTemp       => APUFCMRBDATA_OUT(13),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(13),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(14),
	GlitchData    => APUFCMRBDATA14_GlitchData,
	OutSignalName => "APUFCMRBDATA(14)",
	OutTemp       => APUFCMRBDATA_OUT(14),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(14),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(15),
	GlitchData    => APUFCMRBDATA15_GlitchData,
	OutSignalName => "APUFCMRBDATA(15)",
	OutTemp       => APUFCMRBDATA_OUT(15),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(15),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(16),
	GlitchData    => APUFCMRBDATA16_GlitchData,
	OutSignalName => "APUFCMRBDATA(16)",
	OutTemp       => APUFCMRBDATA_OUT(16),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(16),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(17),
	GlitchData    => APUFCMRBDATA17_GlitchData,
	OutSignalName => "APUFCMRBDATA(17)",
	OutTemp       => APUFCMRBDATA_OUT(17),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(17),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(18),
	GlitchData    => APUFCMRBDATA18_GlitchData,
	OutSignalName => "APUFCMRBDATA(18)",
	OutTemp       => APUFCMRBDATA_OUT(18),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(18),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(19),
	GlitchData    => APUFCMRBDATA19_GlitchData,
	OutSignalName => "APUFCMRBDATA(19)",
	OutTemp       => APUFCMRBDATA_OUT(19),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(19),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(20),
	GlitchData    => APUFCMRBDATA20_GlitchData,
	OutSignalName => "APUFCMRBDATA(20)",
	OutTemp       => APUFCMRBDATA_OUT(20),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(20),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(21),
	GlitchData    => APUFCMRBDATA21_GlitchData,
	OutSignalName => "APUFCMRBDATA(21)",
	OutTemp       => APUFCMRBDATA_OUT(21),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(21),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(22),
	GlitchData    => APUFCMRBDATA22_GlitchData,
	OutSignalName => "APUFCMRBDATA(22)",
	OutTemp       => APUFCMRBDATA_OUT(22),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(22),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(23),
	GlitchData    => APUFCMRBDATA23_GlitchData,
	OutSignalName => "APUFCMRBDATA(23)",
	OutTemp       => APUFCMRBDATA_OUT(23),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(23),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(24),
	GlitchData    => APUFCMRBDATA24_GlitchData,
	OutSignalName => "APUFCMRBDATA(24)",
	OutTemp       => APUFCMRBDATA_OUT(24),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(24),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(25),
	GlitchData    => APUFCMRBDATA25_GlitchData,
	OutSignalName => "APUFCMRBDATA(25)",
	OutTemp       => APUFCMRBDATA_OUT(25),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(25),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(26),
	GlitchData    => APUFCMRBDATA26_GlitchData,
	OutSignalName => "APUFCMRBDATA(26)",
	OutTemp       => APUFCMRBDATA_OUT(26),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(26),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(27),
	GlitchData    => APUFCMRBDATA27_GlitchData,
	OutSignalName => "APUFCMRBDATA(27)",
	OutTemp       => APUFCMRBDATA_OUT(27),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(27),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(28),
	GlitchData    => APUFCMRBDATA28_GlitchData,
	OutSignalName => "APUFCMRBDATA(28)",
	OutTemp       => APUFCMRBDATA_OUT(28),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(28),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(29),
	GlitchData    => APUFCMRBDATA29_GlitchData,
	OutSignalName => "APUFCMRBDATA(29)",
	OutTemp       => APUFCMRBDATA_OUT(29),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(29),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(30),
	GlitchData    => APUFCMRBDATA30_GlitchData,
	OutSignalName => "APUFCMRBDATA(30)",
	OutTemp       => APUFCMRBDATA_OUT(30),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(30),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMRBDATA(31),
	GlitchData    => APUFCMRBDATA31_GlitchData,
	OutSignalName => "APUFCMRBDATA(31)",
	OutTemp       => APUFCMRBDATA_OUT(31),
	Paths       => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMRBDATA(31),TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMRBDATA(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => APUFCMWRITEBACKOK,
	GlitchData    => APUFCMWRITEBACKOK_GlitchData,
	OutSignalName => "APUFCMWRITEBACKOK",
	OutTemp       => APUFCMWRITEBACKOK_OUT,
	Paths         => (0 => (CPMFCMCLK_dly'last_event, tpd_CPMFCMCLK_APUFCMWRITEBACKOK,TRUE)),
	 DefaultDelay =>  tpd_CPMFCMCLK_APUFCMWRITEBACKOK, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440CPMCORESLEEPREQ,
	GlitchData    => C440CPMCORESLEEPREQ_GlitchData,
	OutSignalName => "C440CPMCORESLEEPREQ",
	OutTemp       => C440CPMCORESLEEPREQ_OUT,
	Paths         => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440CPMCORESLEEPREQ,TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440CPMCORESLEEPREQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440CPMDECIRPTREQ,
	GlitchData    => C440CPMDECIRPTREQ_GlitchData,
	OutSignalName => "C440CPMDECIRPTREQ",
	OutTemp       => C440CPMDECIRPTREQ_OUT,
	Paths         => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440CPMDECIRPTREQ,TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440CPMDECIRPTREQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440CPMFITIRPTREQ,
	GlitchData    => C440CPMFITIRPTREQ_GlitchData,
	OutSignalName => "C440CPMFITIRPTREQ",
	OutTemp       => C440CPMFITIRPTREQ_OUT,
	Paths         => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440CPMFITIRPTREQ,TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440CPMFITIRPTREQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440CPMMSRCE,
	GlitchData    => C440CPMMSRCE_GlitchData,
	OutSignalName => "C440CPMMSRCE",
	OutTemp       => C440CPMMSRCE_OUT,
	Paths         => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440CPMMSRCE,TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440CPMMSRCE, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440CPMMSREE,
	GlitchData    => C440CPMMSREE_GlitchData,
	OutSignalName => "C440CPMMSREE",
	OutTemp       => C440CPMMSREE_OUT,
	Paths         => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440CPMMSREE,TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440CPMMSREE, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440CPMTIMERRESETREQ,
	GlitchData    => C440CPMTIMERRESETREQ_GlitchData,
	OutSignalName => "C440CPMTIMERRESETREQ",
	OutTemp       => C440CPMTIMERRESETREQ_OUT,
	Paths         => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440CPMTIMERRESETREQ,TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440CPMTIMERRESETREQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440CPMWDIRPTREQ,
	GlitchData    => C440CPMWDIRPTREQ_GlitchData,
	OutSignalName => "C440CPMWDIRPTREQ",
	OutTemp       => C440CPMWDIRPTREQ_OUT,
	Paths         => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440CPMWDIRPTREQ,TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440CPMWDIRPTREQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(0),
	GlitchData    => C440DBGSYSTEMCONTROL0_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(0)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(0),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(0),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(1),
	GlitchData    => C440DBGSYSTEMCONTROL1_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(1)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(1),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(1),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(2),
	GlitchData    => C440DBGSYSTEMCONTROL2_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(2)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(2),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(2),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(3),
	GlitchData    => C440DBGSYSTEMCONTROL3_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(3)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(3),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(3),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(4),
	GlitchData    => C440DBGSYSTEMCONTROL4_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(4)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(4),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(4),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(5),
	GlitchData    => C440DBGSYSTEMCONTROL5_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(5)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(5),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(5),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(6),
	GlitchData    => C440DBGSYSTEMCONTROL6_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(6)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(6),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(6),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440DBGSYSTEMCONTROL(7),
	GlitchData    => C440DBGSYSTEMCONTROL7_GlitchData,
	OutSignalName => "C440DBGSYSTEMCONTROL(7)",
	OutTemp       => C440DBGSYSTEMCONTROL_OUT(7),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(7),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440DBGSYSTEMCONTROL(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440JTGTDO,
	GlitchData    => C440JTGTDO_GlitchData,
	OutSignalName => "C440JTGTDO",
	OutTemp       => C440JTGTDO_OUT,
	Paths         => (0 => (JTGC440TCK_dly'last_event, tpd_JTGC440TCK_C440JTGTDO,TRUE)),
	 DefaultDelay =>  tpd_JTGC440TCK_C440JTGTDO, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440JTGTDOEN,
	GlitchData    => C440JTGTDOEN_GlitchData,
	OutSignalName => "C440JTGTDOEN",
	OutTemp       => C440JTGTDOEN_OUT,
	Paths         => (0 => (JTGC440TCK_dly'last_event, tpd_JTGC440TCK_C440JTGTDOEN,TRUE)),
	 DefaultDelay =>  tpd_JTGC440TCK_C440JTGTDOEN, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440MACHINECHECK,
	GlitchData    => C440MACHINECHECK_GlitchData,
	OutSignalName => "C440MACHINECHECK",
	OutTemp       => C440MACHINECHECK_OUT,
	Paths         => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440MACHINECHECK,TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440MACHINECHECK, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440RSTCHIPRESETREQ,
	GlitchData    => C440RSTCHIPRESETREQ_GlitchData,
	OutSignalName => "C440RSTCHIPRESETREQ",
	OutTemp       => C440RSTCHIPRESETREQ_OUT,
	Paths         => (0 => (CPMINTERCONNECTCLK_dly'last_event, tpd_CPMINTERCONNECTCLK_C440RSTCHIPRESETREQ,TRUE)),
	 DefaultDelay =>  tpd_CPMINTERCONNECTCLK_C440RSTCHIPRESETREQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440RSTCORERESETREQ,
	GlitchData    => C440RSTCORERESETREQ_GlitchData,
	OutSignalName => "C440RSTCORERESETREQ",
	OutTemp       => C440RSTCORERESETREQ_OUT,
	Paths         => (0 => (CPMINTERCONNECTCLK_dly'last_event, tpd_CPMINTERCONNECTCLK_C440RSTCORERESETREQ,TRUE)),
	 DefaultDelay =>  tpd_CPMINTERCONNECTCLK_C440RSTCORERESETREQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440RSTSYSTEMRESETREQ,
	GlitchData    => C440RSTSYSTEMRESETREQ_GlitchData,
	OutSignalName => "C440RSTSYSTEMRESETREQ",
	OutTemp       => C440RSTSYSTEMRESETREQ_OUT,
	Paths         => (0 => (CPMINTERCONNECTCLK_dly'last_event, tpd_CPMINTERCONNECTCLK_C440RSTSYSTEMRESETREQ,TRUE)),
	 DefaultDelay =>  tpd_CPMINTERCONNECTCLK_C440RSTSYSTEMRESETREQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCBRANCHSTATUS(0),
	GlitchData    => C440TRCBRANCHSTATUS0_GlitchData,
	OutSignalName => "C440TRCBRANCHSTATUS(0)",
	OutTemp       => C440TRCBRANCHSTATUS_OUT(0),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCBRANCHSTATUS(0),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCBRANCHSTATUS(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCBRANCHSTATUS(1),
	GlitchData    => C440TRCBRANCHSTATUS1_GlitchData,
	OutSignalName => "C440TRCBRANCHSTATUS(1)",
	OutTemp       => C440TRCBRANCHSTATUS_OUT(1),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCBRANCHSTATUS(1),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCBRANCHSTATUS(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCBRANCHSTATUS(2),
	GlitchData    => C440TRCBRANCHSTATUS2_GlitchData,
	OutSignalName => "C440TRCBRANCHSTATUS(2)",
	OutTemp       => C440TRCBRANCHSTATUS_OUT(2),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCBRANCHSTATUS(2),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCBRANCHSTATUS(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCCYCLE,
	GlitchData    => C440TRCCYCLE_GlitchData,
	OutSignalName => "C440TRCCYCLE",
	OutTemp       => C440TRCCYCLE_OUT,
	Paths         => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCCYCLE,TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCCYCLE, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCEXECUTIONSTATUS(0),
	GlitchData    => C440TRCEXECUTIONSTATUS0_GlitchData,
	OutSignalName => "C440TRCEXECUTIONSTATUS(0)",
	OutTemp       => C440TRCEXECUTIONSTATUS_OUT(0),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCEXECUTIONSTATUS(0),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCEXECUTIONSTATUS(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCEXECUTIONSTATUS(1),
	GlitchData    => C440TRCEXECUTIONSTATUS1_GlitchData,
	OutSignalName => "C440TRCEXECUTIONSTATUS(1)",
	OutTemp       => C440TRCEXECUTIONSTATUS_OUT(1),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCEXECUTIONSTATUS(1),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCEXECUTIONSTATUS(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCEXECUTIONSTATUS(2),
	GlitchData    => C440TRCEXECUTIONSTATUS2_GlitchData,
	OutSignalName => "C440TRCEXECUTIONSTATUS(2)",
	OutTemp       => C440TRCEXECUTIONSTATUS_OUT(2),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCEXECUTIONSTATUS(2),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCEXECUTIONSTATUS(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCEXECUTIONSTATUS(3),
	GlitchData    => C440TRCEXECUTIONSTATUS3_GlitchData,
	OutSignalName => "C440TRCEXECUTIONSTATUS(3)",
	OutTemp       => C440TRCEXECUTIONSTATUS_OUT(3),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCEXECUTIONSTATUS(3),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCEXECUTIONSTATUS(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCEXECUTIONSTATUS(4),
	GlitchData    => C440TRCEXECUTIONSTATUS4_GlitchData,
	OutSignalName => "C440TRCEXECUTIONSTATUS(4)",
	OutTemp       => C440TRCEXECUTIONSTATUS_OUT(4),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCEXECUTIONSTATUS(4),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCEXECUTIONSTATUS(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRACESTATUS(0),
	GlitchData    => C440TRCTRACESTATUS0_GlitchData,
	OutSignalName => "C440TRCTRACESTATUS(0)",
	OutTemp       => C440TRCTRACESTATUS_OUT(0),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRACESTATUS(0),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRACESTATUS(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRACESTATUS(1),
	GlitchData    => C440TRCTRACESTATUS1_GlitchData,
	OutSignalName => "C440TRCTRACESTATUS(1)",
	OutTemp       => C440TRCTRACESTATUS_OUT(1),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRACESTATUS(1),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRACESTATUS(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRACESTATUS(2),
	GlitchData    => C440TRCTRACESTATUS2_GlitchData,
	OutSignalName => "C440TRCTRACESTATUS(2)",
	OutTemp       => C440TRCTRACESTATUS_OUT(2),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRACESTATUS(2),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRACESTATUS(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRACESTATUS(3),
	GlitchData    => C440TRCTRACESTATUS3_GlitchData,
	OutSignalName => "C440TRCTRACESTATUS(3)",
	OutTemp       => C440TRCTRACESTATUS_OUT(3),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRACESTATUS(3),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRACESTATUS(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRACESTATUS(4),
	GlitchData    => C440TRCTRACESTATUS4_GlitchData,
	OutSignalName => "C440TRCTRACESTATUS(4)",
	OutTemp       => C440TRCTRACESTATUS_OUT(4),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRACESTATUS(4),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRACESTATUS(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRACESTATUS(5),
	GlitchData    => C440TRCTRACESTATUS5_GlitchData,
	OutSignalName => "C440TRCTRACESTATUS(5)",
	OutTemp       => C440TRCTRACESTATUS_OUT(5),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRACESTATUS(5),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRACESTATUS(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRACESTATUS(6),
	GlitchData    => C440TRCTRACESTATUS6_GlitchData,
	OutSignalName => "C440TRCTRACESTATUS(6)",
	OutTemp       => C440TRCTRACESTATUS_OUT(6),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRACESTATUS(6),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRACESTATUS(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTOUT,
	GlitchData    => C440TRCTRIGGEREVENTOUT_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTOUT",
	OutTemp       => C440TRCTRIGGEREVENTOUT_OUT,
	Paths         => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTOUT,TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTOUT, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(0),
	GlitchData    => C440TRCTRIGGEREVENTTYPE0_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(0)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(0),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(0),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(1),
	GlitchData    => C440TRCTRIGGEREVENTTYPE1_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(1)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(1),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(1),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(2),
	GlitchData    => C440TRCTRIGGEREVENTTYPE2_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(2)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(2),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(2),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(3),
	GlitchData    => C440TRCTRIGGEREVENTTYPE3_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(3)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(3),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(3),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(4),
	GlitchData    => C440TRCTRIGGEREVENTTYPE4_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(4)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(4),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(4),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(5),
	GlitchData    => C440TRCTRIGGEREVENTTYPE5_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(5)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(5),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(5),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(6),
	GlitchData    => C440TRCTRIGGEREVENTTYPE6_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(6)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(6),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(6),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(7),
	GlitchData    => C440TRCTRIGGEREVENTTYPE7_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(7)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(7),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(7),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(8),
	GlitchData    => C440TRCTRIGGEREVENTTYPE8_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(8)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(8),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(8),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(9),
	GlitchData    => C440TRCTRIGGEREVENTTYPE9_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(9)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(9),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(9),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(10),
	GlitchData    => C440TRCTRIGGEREVENTTYPE10_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(10)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(10),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(10),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(11),
	GlitchData    => C440TRCTRIGGEREVENTTYPE11_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(11)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(11),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(11),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(12),
	GlitchData    => C440TRCTRIGGEREVENTTYPE12_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(12)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(12),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(12),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => C440TRCTRIGGEREVENTTYPE(13),
	GlitchData    => C440TRCTRIGGEREVENTTYPE13_GlitchData,
	OutSignalName => "C440TRCTRIGGEREVENTTYPE(13)",
	OutTemp       => C440TRCTRIGGEREVENTTYPE_OUT(13),
	Paths       => (0 => (CPMC440CLK_dly'last_event, tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(13),TRUE)),
	 DefaultDelay =>  tpd_CPMC440CLK_C440TRCTRIGGEREVENTTYPE(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(0),
	GlitchData    => MIMCADDRESS0_GlitchData,
	OutSignalName => "MIMCADDRESS(0)",
	OutTemp       => MIMCADDRESS_OUT(0),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(0),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(1),
	GlitchData    => MIMCADDRESS1_GlitchData,
	OutSignalName => "MIMCADDRESS(1)",
	OutTemp       => MIMCADDRESS_OUT(1),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(1),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(2),
	GlitchData    => MIMCADDRESS2_GlitchData,
	OutSignalName => "MIMCADDRESS(2)",
	OutTemp       => MIMCADDRESS_OUT(2),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(2),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(3),
	GlitchData    => MIMCADDRESS3_GlitchData,
	OutSignalName => "MIMCADDRESS(3)",
	OutTemp       => MIMCADDRESS_OUT(3),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(3),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(4),
	GlitchData    => MIMCADDRESS4_GlitchData,
	OutSignalName => "MIMCADDRESS(4)",
	OutTemp       => MIMCADDRESS_OUT(4),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(4),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(5),
	GlitchData    => MIMCADDRESS5_GlitchData,
	OutSignalName => "MIMCADDRESS(5)",
	OutTemp       => MIMCADDRESS_OUT(5),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(5),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(6),
	GlitchData    => MIMCADDRESS6_GlitchData,
	OutSignalName => "MIMCADDRESS(6)",
	OutTemp       => MIMCADDRESS_OUT(6),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(6),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(7),
	GlitchData    => MIMCADDRESS7_GlitchData,
	OutSignalName => "MIMCADDRESS(7)",
	OutTemp       => MIMCADDRESS_OUT(7),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(7),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(8),
	GlitchData    => MIMCADDRESS8_GlitchData,
	OutSignalName => "MIMCADDRESS(8)",
	OutTemp       => MIMCADDRESS_OUT(8),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(8),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(9),
	GlitchData    => MIMCADDRESS9_GlitchData,
	OutSignalName => "MIMCADDRESS(9)",
	OutTemp       => MIMCADDRESS_OUT(9),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(9),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(10),
	GlitchData    => MIMCADDRESS10_GlitchData,
	OutSignalName => "MIMCADDRESS(10)",
	OutTemp       => MIMCADDRESS_OUT(10),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(10),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(11),
	GlitchData    => MIMCADDRESS11_GlitchData,
	OutSignalName => "MIMCADDRESS(11)",
	OutTemp       => MIMCADDRESS_OUT(11),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(11),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(12),
	GlitchData    => MIMCADDRESS12_GlitchData,
	OutSignalName => "MIMCADDRESS(12)",
	OutTemp       => MIMCADDRESS_OUT(12),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(12),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(13),
	GlitchData    => MIMCADDRESS13_GlitchData,
	OutSignalName => "MIMCADDRESS(13)",
	OutTemp       => MIMCADDRESS_OUT(13),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(13),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(14),
	GlitchData    => MIMCADDRESS14_GlitchData,
	OutSignalName => "MIMCADDRESS(14)",
	OutTemp       => MIMCADDRESS_OUT(14),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(14),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(15),
	GlitchData    => MIMCADDRESS15_GlitchData,
	OutSignalName => "MIMCADDRESS(15)",
	OutTemp       => MIMCADDRESS_OUT(15),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(15),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(16),
	GlitchData    => MIMCADDRESS16_GlitchData,
	OutSignalName => "MIMCADDRESS(16)",
	OutTemp       => MIMCADDRESS_OUT(16),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(16),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(17),
	GlitchData    => MIMCADDRESS17_GlitchData,
	OutSignalName => "MIMCADDRESS(17)",
	OutTemp       => MIMCADDRESS_OUT(17),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(17),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(18),
	GlitchData    => MIMCADDRESS18_GlitchData,
	OutSignalName => "MIMCADDRESS(18)",
	OutTemp       => MIMCADDRESS_OUT(18),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(18),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(19),
	GlitchData    => MIMCADDRESS19_GlitchData,
	OutSignalName => "MIMCADDRESS(19)",
	OutTemp       => MIMCADDRESS_OUT(19),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(19),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(20),
	GlitchData    => MIMCADDRESS20_GlitchData,
	OutSignalName => "MIMCADDRESS(20)",
	OutTemp       => MIMCADDRESS_OUT(20),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(20),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(21),
	GlitchData    => MIMCADDRESS21_GlitchData,
	OutSignalName => "MIMCADDRESS(21)",
	OutTemp       => MIMCADDRESS_OUT(21),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(21),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(22),
	GlitchData    => MIMCADDRESS22_GlitchData,
	OutSignalName => "MIMCADDRESS(22)",
	OutTemp       => MIMCADDRESS_OUT(22),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(22),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(23),
	GlitchData    => MIMCADDRESS23_GlitchData,
	OutSignalName => "MIMCADDRESS(23)",
	OutTemp       => MIMCADDRESS_OUT(23),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(23),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(24),
	GlitchData    => MIMCADDRESS24_GlitchData,
	OutSignalName => "MIMCADDRESS(24)",
	OutTemp       => MIMCADDRESS_OUT(24),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(24),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(25),
	GlitchData    => MIMCADDRESS25_GlitchData,
	OutSignalName => "MIMCADDRESS(25)",
	OutTemp       => MIMCADDRESS_OUT(25),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(25),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(26),
	GlitchData    => MIMCADDRESS26_GlitchData,
	OutSignalName => "MIMCADDRESS(26)",
	OutTemp       => MIMCADDRESS_OUT(26),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(26),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(27),
	GlitchData    => MIMCADDRESS27_GlitchData,
	OutSignalName => "MIMCADDRESS(27)",
	OutTemp       => MIMCADDRESS_OUT(27),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(27),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(28),
	GlitchData    => MIMCADDRESS28_GlitchData,
	OutSignalName => "MIMCADDRESS(28)",
	OutTemp       => MIMCADDRESS_OUT(28),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(28),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(29),
	GlitchData    => MIMCADDRESS29_GlitchData,
	OutSignalName => "MIMCADDRESS(29)",
	OutTemp       => MIMCADDRESS_OUT(29),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(29),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(30),
	GlitchData    => MIMCADDRESS30_GlitchData,
	OutSignalName => "MIMCADDRESS(30)",
	OutTemp       => MIMCADDRESS_OUT(30),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(30),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(31),
	GlitchData    => MIMCADDRESS31_GlitchData,
	OutSignalName => "MIMCADDRESS(31)",
	OutTemp       => MIMCADDRESS_OUT(31),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(31),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(32),
	GlitchData    => MIMCADDRESS32_GlitchData,
	OutSignalName => "MIMCADDRESS(32)",
	OutTemp       => MIMCADDRESS_OUT(32),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(32),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(32), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(33),
	GlitchData    => MIMCADDRESS33_GlitchData,
	OutSignalName => "MIMCADDRESS(33)",
	OutTemp       => MIMCADDRESS_OUT(33),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(33),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(33), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(34),
	GlitchData    => MIMCADDRESS34_GlitchData,
	OutSignalName => "MIMCADDRESS(34)",
	OutTemp       => MIMCADDRESS_OUT(34),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(34),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(34), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESS(35),
	GlitchData    => MIMCADDRESS35_GlitchData,
	OutSignalName => "MIMCADDRESS(35)",
	OutTemp       => MIMCADDRESS_OUT(35),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESS(35),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESS(35), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCADDRESSVALID,
	GlitchData    => MIMCADDRESSVALID_GlitchData,
	OutSignalName => "MIMCADDRESSVALID",
	OutTemp       => MIMCADDRESSVALID_OUT,
	Paths         => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCADDRESSVALID,TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCADDRESSVALID, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBANKCONFLICT,
	GlitchData    => MIMCBANKCONFLICT_GlitchData,
	OutSignalName => "MIMCBANKCONFLICT",
	OutTemp       => MIMCBANKCONFLICT_OUT,
	Paths         => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBANKCONFLICT,TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBANKCONFLICT, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(0),
	GlitchData    => MIMCBYTEENABLE0_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(0)",
	OutTemp       => MIMCBYTEENABLE_OUT(0),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(0),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(1),
	GlitchData    => MIMCBYTEENABLE1_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(1)",
	OutTemp       => MIMCBYTEENABLE_OUT(1),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(1),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(2),
	GlitchData    => MIMCBYTEENABLE2_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(2)",
	OutTemp       => MIMCBYTEENABLE_OUT(2),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(2),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(3),
	GlitchData    => MIMCBYTEENABLE3_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(3)",
	OutTemp       => MIMCBYTEENABLE_OUT(3),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(3),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(4),
	GlitchData    => MIMCBYTEENABLE4_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(4)",
	OutTemp       => MIMCBYTEENABLE_OUT(4),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(4),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(5),
	GlitchData    => MIMCBYTEENABLE5_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(5)",
	OutTemp       => MIMCBYTEENABLE_OUT(5),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(5),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(6),
	GlitchData    => MIMCBYTEENABLE6_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(6)",
	OutTemp       => MIMCBYTEENABLE_OUT(6),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(6),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(7),
	GlitchData    => MIMCBYTEENABLE7_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(7)",
	OutTemp       => MIMCBYTEENABLE_OUT(7),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(7),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(8),
	GlitchData    => MIMCBYTEENABLE8_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(8)",
	OutTemp       => MIMCBYTEENABLE_OUT(8),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(8),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(9),
	GlitchData    => MIMCBYTEENABLE9_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(9)",
	OutTemp       => MIMCBYTEENABLE_OUT(9),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(9),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(10),
	GlitchData    => MIMCBYTEENABLE10_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(10)",
	OutTemp       => MIMCBYTEENABLE_OUT(10),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(10),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(11),
	GlitchData    => MIMCBYTEENABLE11_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(11)",
	OutTemp       => MIMCBYTEENABLE_OUT(11),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(11),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(12),
	GlitchData    => MIMCBYTEENABLE12_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(12)",
	OutTemp       => MIMCBYTEENABLE_OUT(12),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(12),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(13),
	GlitchData    => MIMCBYTEENABLE13_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(13)",
	OutTemp       => MIMCBYTEENABLE_OUT(13),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(13),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(14),
	GlitchData    => MIMCBYTEENABLE14_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(14)",
	OutTemp       => MIMCBYTEENABLE_OUT(14),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(14),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCBYTEENABLE(15),
	GlitchData    => MIMCBYTEENABLE15_GlitchData,
	OutSignalName => "MIMCBYTEENABLE(15)",
	OutTemp       => MIMCBYTEENABLE_OUT(15),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCBYTEENABLE(15),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCBYTEENABLE(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCREADNOTWRITE,
	GlitchData    => MIMCREADNOTWRITE_GlitchData,
	OutSignalName => "MIMCREADNOTWRITE",
	OutTemp       => MIMCREADNOTWRITE_OUT,
	Paths         => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCREADNOTWRITE,TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCREADNOTWRITE, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCROWCONFLICT,
	GlitchData    => MIMCROWCONFLICT_GlitchData,
	OutSignalName => "MIMCROWCONFLICT",
	OutTemp       => MIMCROWCONFLICT_OUT,
	Paths         => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCROWCONFLICT,TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCROWCONFLICT, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(0),
	GlitchData    => MIMCWRITEDATA0_GlitchData,
	OutSignalName => "MIMCWRITEDATA(0)",
	OutTemp       => MIMCWRITEDATA_OUT(0),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(0),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(1),
	GlitchData    => MIMCWRITEDATA1_GlitchData,
	OutSignalName => "MIMCWRITEDATA(1)",
	OutTemp       => MIMCWRITEDATA_OUT(1),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(1),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(2),
	GlitchData    => MIMCWRITEDATA2_GlitchData,
	OutSignalName => "MIMCWRITEDATA(2)",
	OutTemp       => MIMCWRITEDATA_OUT(2),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(2),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(3),
	GlitchData    => MIMCWRITEDATA3_GlitchData,
	OutSignalName => "MIMCWRITEDATA(3)",
	OutTemp       => MIMCWRITEDATA_OUT(3),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(3),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(4),
	GlitchData    => MIMCWRITEDATA4_GlitchData,
	OutSignalName => "MIMCWRITEDATA(4)",
	OutTemp       => MIMCWRITEDATA_OUT(4),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(4),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(5),
	GlitchData    => MIMCWRITEDATA5_GlitchData,
	OutSignalName => "MIMCWRITEDATA(5)",
	OutTemp       => MIMCWRITEDATA_OUT(5),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(5),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(6),
	GlitchData    => MIMCWRITEDATA6_GlitchData,
	OutSignalName => "MIMCWRITEDATA(6)",
	OutTemp       => MIMCWRITEDATA_OUT(6),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(6),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(7),
	GlitchData    => MIMCWRITEDATA7_GlitchData,
	OutSignalName => "MIMCWRITEDATA(7)",
	OutTemp       => MIMCWRITEDATA_OUT(7),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(7),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(8),
	GlitchData    => MIMCWRITEDATA8_GlitchData,
	OutSignalName => "MIMCWRITEDATA(8)",
	OutTemp       => MIMCWRITEDATA_OUT(8),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(8),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(9),
	GlitchData    => MIMCWRITEDATA9_GlitchData,
	OutSignalName => "MIMCWRITEDATA(9)",
	OutTemp       => MIMCWRITEDATA_OUT(9),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(9),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(10),
	GlitchData    => MIMCWRITEDATA10_GlitchData,
	OutSignalName => "MIMCWRITEDATA(10)",
	OutTemp       => MIMCWRITEDATA_OUT(10),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(10),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(11),
	GlitchData    => MIMCWRITEDATA11_GlitchData,
	OutSignalName => "MIMCWRITEDATA(11)",
	OutTemp       => MIMCWRITEDATA_OUT(11),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(11),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(12),
	GlitchData    => MIMCWRITEDATA12_GlitchData,
	OutSignalName => "MIMCWRITEDATA(12)",
	OutTemp       => MIMCWRITEDATA_OUT(12),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(12),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(13),
	GlitchData    => MIMCWRITEDATA13_GlitchData,
	OutSignalName => "MIMCWRITEDATA(13)",
	OutTemp       => MIMCWRITEDATA_OUT(13),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(13),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(14),
	GlitchData    => MIMCWRITEDATA14_GlitchData,
	OutSignalName => "MIMCWRITEDATA(14)",
	OutTemp       => MIMCWRITEDATA_OUT(14),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(14),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(15),
	GlitchData    => MIMCWRITEDATA15_GlitchData,
	OutSignalName => "MIMCWRITEDATA(15)",
	OutTemp       => MIMCWRITEDATA_OUT(15),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(15),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(16),
	GlitchData    => MIMCWRITEDATA16_GlitchData,
	OutSignalName => "MIMCWRITEDATA(16)",
	OutTemp       => MIMCWRITEDATA_OUT(16),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(16),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(17),
	GlitchData    => MIMCWRITEDATA17_GlitchData,
	OutSignalName => "MIMCWRITEDATA(17)",
	OutTemp       => MIMCWRITEDATA_OUT(17),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(17),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(18),
	GlitchData    => MIMCWRITEDATA18_GlitchData,
	OutSignalName => "MIMCWRITEDATA(18)",
	OutTemp       => MIMCWRITEDATA_OUT(18),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(18),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(19),
	GlitchData    => MIMCWRITEDATA19_GlitchData,
	OutSignalName => "MIMCWRITEDATA(19)",
	OutTemp       => MIMCWRITEDATA_OUT(19),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(19),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(20),
	GlitchData    => MIMCWRITEDATA20_GlitchData,
	OutSignalName => "MIMCWRITEDATA(20)",
	OutTemp       => MIMCWRITEDATA_OUT(20),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(20),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(21),
	GlitchData    => MIMCWRITEDATA21_GlitchData,
	OutSignalName => "MIMCWRITEDATA(21)",
	OutTemp       => MIMCWRITEDATA_OUT(21),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(21),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(22),
	GlitchData    => MIMCWRITEDATA22_GlitchData,
	OutSignalName => "MIMCWRITEDATA(22)",
	OutTemp       => MIMCWRITEDATA_OUT(22),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(22),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(23),
	GlitchData    => MIMCWRITEDATA23_GlitchData,
	OutSignalName => "MIMCWRITEDATA(23)",
	OutTemp       => MIMCWRITEDATA_OUT(23),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(23),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(24),
	GlitchData    => MIMCWRITEDATA24_GlitchData,
	OutSignalName => "MIMCWRITEDATA(24)",
	OutTemp       => MIMCWRITEDATA_OUT(24),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(24),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(25),
	GlitchData    => MIMCWRITEDATA25_GlitchData,
	OutSignalName => "MIMCWRITEDATA(25)",
	OutTemp       => MIMCWRITEDATA_OUT(25),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(25),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(26),
	GlitchData    => MIMCWRITEDATA26_GlitchData,
	OutSignalName => "MIMCWRITEDATA(26)",
	OutTemp       => MIMCWRITEDATA_OUT(26),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(26),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(27),
	GlitchData    => MIMCWRITEDATA27_GlitchData,
	OutSignalName => "MIMCWRITEDATA(27)",
	OutTemp       => MIMCWRITEDATA_OUT(27),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(27),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(28),
	GlitchData    => MIMCWRITEDATA28_GlitchData,
	OutSignalName => "MIMCWRITEDATA(28)",
	OutTemp       => MIMCWRITEDATA_OUT(28),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(28),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(29),
	GlitchData    => MIMCWRITEDATA29_GlitchData,
	OutSignalName => "MIMCWRITEDATA(29)",
	OutTemp       => MIMCWRITEDATA_OUT(29),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(29),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(30),
	GlitchData    => MIMCWRITEDATA30_GlitchData,
	OutSignalName => "MIMCWRITEDATA(30)",
	OutTemp       => MIMCWRITEDATA_OUT(30),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(30),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(31),
	GlitchData    => MIMCWRITEDATA31_GlitchData,
	OutSignalName => "MIMCWRITEDATA(31)",
	OutTemp       => MIMCWRITEDATA_OUT(31),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(31),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(32),
	GlitchData    => MIMCWRITEDATA32_GlitchData,
	OutSignalName => "MIMCWRITEDATA(32)",
	OutTemp       => MIMCWRITEDATA_OUT(32),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(32),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(32), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(33),
	GlitchData    => MIMCWRITEDATA33_GlitchData,
	OutSignalName => "MIMCWRITEDATA(33)",
	OutTemp       => MIMCWRITEDATA_OUT(33),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(33),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(33), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(34),
	GlitchData    => MIMCWRITEDATA34_GlitchData,
	OutSignalName => "MIMCWRITEDATA(34)",
	OutTemp       => MIMCWRITEDATA_OUT(34),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(34),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(34), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(35),
	GlitchData    => MIMCWRITEDATA35_GlitchData,
	OutSignalName => "MIMCWRITEDATA(35)",
	OutTemp       => MIMCWRITEDATA_OUT(35),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(35),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(35), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(36),
	GlitchData    => MIMCWRITEDATA36_GlitchData,
	OutSignalName => "MIMCWRITEDATA(36)",
	OutTemp       => MIMCWRITEDATA_OUT(36),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(36),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(36), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(37),
	GlitchData    => MIMCWRITEDATA37_GlitchData,
	OutSignalName => "MIMCWRITEDATA(37)",
	OutTemp       => MIMCWRITEDATA_OUT(37),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(37),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(37), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(38),
	GlitchData    => MIMCWRITEDATA38_GlitchData,
	OutSignalName => "MIMCWRITEDATA(38)",
	OutTemp       => MIMCWRITEDATA_OUT(38),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(38),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(38), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(39),
	GlitchData    => MIMCWRITEDATA39_GlitchData,
	OutSignalName => "MIMCWRITEDATA(39)",
	OutTemp       => MIMCWRITEDATA_OUT(39),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(39),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(39), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(40),
	GlitchData    => MIMCWRITEDATA40_GlitchData,
	OutSignalName => "MIMCWRITEDATA(40)",
	OutTemp       => MIMCWRITEDATA_OUT(40),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(40),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(40), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(41),
	GlitchData    => MIMCWRITEDATA41_GlitchData,
	OutSignalName => "MIMCWRITEDATA(41)",
	OutTemp       => MIMCWRITEDATA_OUT(41),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(41),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(41), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(42),
	GlitchData    => MIMCWRITEDATA42_GlitchData,
	OutSignalName => "MIMCWRITEDATA(42)",
	OutTemp       => MIMCWRITEDATA_OUT(42),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(42),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(42), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(43),
	GlitchData    => MIMCWRITEDATA43_GlitchData,
	OutSignalName => "MIMCWRITEDATA(43)",
	OutTemp       => MIMCWRITEDATA_OUT(43),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(43),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(43), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(44),
	GlitchData    => MIMCWRITEDATA44_GlitchData,
	OutSignalName => "MIMCWRITEDATA(44)",
	OutTemp       => MIMCWRITEDATA_OUT(44),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(44),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(44), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(45),
	GlitchData    => MIMCWRITEDATA45_GlitchData,
	OutSignalName => "MIMCWRITEDATA(45)",
	OutTemp       => MIMCWRITEDATA_OUT(45),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(45),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(45), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(46),
	GlitchData    => MIMCWRITEDATA46_GlitchData,
	OutSignalName => "MIMCWRITEDATA(46)",
	OutTemp       => MIMCWRITEDATA_OUT(46),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(46),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(46), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(47),
	GlitchData    => MIMCWRITEDATA47_GlitchData,
	OutSignalName => "MIMCWRITEDATA(47)",
	OutTemp       => MIMCWRITEDATA_OUT(47),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(47),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(47), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(48),
	GlitchData    => MIMCWRITEDATA48_GlitchData,
	OutSignalName => "MIMCWRITEDATA(48)",
	OutTemp       => MIMCWRITEDATA_OUT(48),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(48),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(48), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(49),
	GlitchData    => MIMCWRITEDATA49_GlitchData,
	OutSignalName => "MIMCWRITEDATA(49)",
	OutTemp       => MIMCWRITEDATA_OUT(49),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(49),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(49), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(50),
	GlitchData    => MIMCWRITEDATA50_GlitchData,
	OutSignalName => "MIMCWRITEDATA(50)",
	OutTemp       => MIMCWRITEDATA_OUT(50),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(50),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(50), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(51),
	GlitchData    => MIMCWRITEDATA51_GlitchData,
	OutSignalName => "MIMCWRITEDATA(51)",
	OutTemp       => MIMCWRITEDATA_OUT(51),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(51),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(51), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(52),
	GlitchData    => MIMCWRITEDATA52_GlitchData,
	OutSignalName => "MIMCWRITEDATA(52)",
	OutTemp       => MIMCWRITEDATA_OUT(52),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(52),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(52), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(53),
	GlitchData    => MIMCWRITEDATA53_GlitchData,
	OutSignalName => "MIMCWRITEDATA(53)",
	OutTemp       => MIMCWRITEDATA_OUT(53),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(53),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(53), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(54),
	GlitchData    => MIMCWRITEDATA54_GlitchData,
	OutSignalName => "MIMCWRITEDATA(54)",
	OutTemp       => MIMCWRITEDATA_OUT(54),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(54),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(54), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(55),
	GlitchData    => MIMCWRITEDATA55_GlitchData,
	OutSignalName => "MIMCWRITEDATA(55)",
	OutTemp       => MIMCWRITEDATA_OUT(55),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(55),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(55), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(56),
	GlitchData    => MIMCWRITEDATA56_GlitchData,
	OutSignalName => "MIMCWRITEDATA(56)",
	OutTemp       => MIMCWRITEDATA_OUT(56),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(56),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(56), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(57),
	GlitchData    => MIMCWRITEDATA57_GlitchData,
	OutSignalName => "MIMCWRITEDATA(57)",
	OutTemp       => MIMCWRITEDATA_OUT(57),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(57),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(57), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(58),
	GlitchData    => MIMCWRITEDATA58_GlitchData,
	OutSignalName => "MIMCWRITEDATA(58)",
	OutTemp       => MIMCWRITEDATA_OUT(58),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(58),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(58), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(59),
	GlitchData    => MIMCWRITEDATA59_GlitchData,
	OutSignalName => "MIMCWRITEDATA(59)",
	OutTemp       => MIMCWRITEDATA_OUT(59),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(59),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(59), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(60),
	GlitchData    => MIMCWRITEDATA60_GlitchData,
	OutSignalName => "MIMCWRITEDATA(60)",
	OutTemp       => MIMCWRITEDATA_OUT(60),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(60),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(60), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(61),
	GlitchData    => MIMCWRITEDATA61_GlitchData,
	OutSignalName => "MIMCWRITEDATA(61)",
	OutTemp       => MIMCWRITEDATA_OUT(61),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(61),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(61), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(62),
	GlitchData    => MIMCWRITEDATA62_GlitchData,
	OutSignalName => "MIMCWRITEDATA(62)",
	OutTemp       => MIMCWRITEDATA_OUT(62),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(62),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(62), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(63),
	GlitchData    => MIMCWRITEDATA63_GlitchData,
	OutSignalName => "MIMCWRITEDATA(63)",
	OutTemp       => MIMCWRITEDATA_OUT(63),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(63),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(63), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(64),
	GlitchData    => MIMCWRITEDATA64_GlitchData,
	OutSignalName => "MIMCWRITEDATA(64)",
	OutTemp       => MIMCWRITEDATA_OUT(64),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(64),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(64), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(65),
	GlitchData    => MIMCWRITEDATA65_GlitchData,
	OutSignalName => "MIMCWRITEDATA(65)",
	OutTemp       => MIMCWRITEDATA_OUT(65),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(65),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(65), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(66),
	GlitchData    => MIMCWRITEDATA66_GlitchData,
	OutSignalName => "MIMCWRITEDATA(66)",
	OutTemp       => MIMCWRITEDATA_OUT(66),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(66),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(66), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(67),
	GlitchData    => MIMCWRITEDATA67_GlitchData,
	OutSignalName => "MIMCWRITEDATA(67)",
	OutTemp       => MIMCWRITEDATA_OUT(67),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(67),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(67), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(68),
	GlitchData    => MIMCWRITEDATA68_GlitchData,
	OutSignalName => "MIMCWRITEDATA(68)",
	OutTemp       => MIMCWRITEDATA_OUT(68),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(68),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(68), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(69),
	GlitchData    => MIMCWRITEDATA69_GlitchData,
	OutSignalName => "MIMCWRITEDATA(69)",
	OutTemp       => MIMCWRITEDATA_OUT(69),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(69),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(69), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(70),
	GlitchData    => MIMCWRITEDATA70_GlitchData,
	OutSignalName => "MIMCWRITEDATA(70)",
	OutTemp       => MIMCWRITEDATA_OUT(70),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(70),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(70), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(71),
	GlitchData    => MIMCWRITEDATA71_GlitchData,
	OutSignalName => "MIMCWRITEDATA(71)",
	OutTemp       => MIMCWRITEDATA_OUT(71),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(71),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(71), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(72),
	GlitchData    => MIMCWRITEDATA72_GlitchData,
	OutSignalName => "MIMCWRITEDATA(72)",
	OutTemp       => MIMCWRITEDATA_OUT(72),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(72),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(72), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(73),
	GlitchData    => MIMCWRITEDATA73_GlitchData,
	OutSignalName => "MIMCWRITEDATA(73)",
	OutTemp       => MIMCWRITEDATA_OUT(73),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(73),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(73), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(74),
	GlitchData    => MIMCWRITEDATA74_GlitchData,
	OutSignalName => "MIMCWRITEDATA(74)",
	OutTemp       => MIMCWRITEDATA_OUT(74),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(74),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(74), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(75),
	GlitchData    => MIMCWRITEDATA75_GlitchData,
	OutSignalName => "MIMCWRITEDATA(75)",
	OutTemp       => MIMCWRITEDATA_OUT(75),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(75),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(75), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(76),
	GlitchData    => MIMCWRITEDATA76_GlitchData,
	OutSignalName => "MIMCWRITEDATA(76)",
	OutTemp       => MIMCWRITEDATA_OUT(76),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(76),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(76), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(77),
	GlitchData    => MIMCWRITEDATA77_GlitchData,
	OutSignalName => "MIMCWRITEDATA(77)",
	OutTemp       => MIMCWRITEDATA_OUT(77),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(77),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(77), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(78),
	GlitchData    => MIMCWRITEDATA78_GlitchData,
	OutSignalName => "MIMCWRITEDATA(78)",
	OutTemp       => MIMCWRITEDATA_OUT(78),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(78),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(78), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(79),
	GlitchData    => MIMCWRITEDATA79_GlitchData,
	OutSignalName => "MIMCWRITEDATA(79)",
	OutTemp       => MIMCWRITEDATA_OUT(79),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(79),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(79), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(80),
	GlitchData    => MIMCWRITEDATA80_GlitchData,
	OutSignalName => "MIMCWRITEDATA(80)",
	OutTemp       => MIMCWRITEDATA_OUT(80),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(80),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(80), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(81),
	GlitchData    => MIMCWRITEDATA81_GlitchData,
	OutSignalName => "MIMCWRITEDATA(81)",
	OutTemp       => MIMCWRITEDATA_OUT(81),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(81),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(81), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(82),
	GlitchData    => MIMCWRITEDATA82_GlitchData,
	OutSignalName => "MIMCWRITEDATA(82)",
	OutTemp       => MIMCWRITEDATA_OUT(82),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(82),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(82), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(83),
	GlitchData    => MIMCWRITEDATA83_GlitchData,
	OutSignalName => "MIMCWRITEDATA(83)",
	OutTemp       => MIMCWRITEDATA_OUT(83),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(83),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(83), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(84),
	GlitchData    => MIMCWRITEDATA84_GlitchData,
	OutSignalName => "MIMCWRITEDATA(84)",
	OutTemp       => MIMCWRITEDATA_OUT(84),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(84),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(84), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(85),
	GlitchData    => MIMCWRITEDATA85_GlitchData,
	OutSignalName => "MIMCWRITEDATA(85)",
	OutTemp       => MIMCWRITEDATA_OUT(85),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(85),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(85), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(86),
	GlitchData    => MIMCWRITEDATA86_GlitchData,
	OutSignalName => "MIMCWRITEDATA(86)",
	OutTemp       => MIMCWRITEDATA_OUT(86),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(86),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(86), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(87),
	GlitchData    => MIMCWRITEDATA87_GlitchData,
	OutSignalName => "MIMCWRITEDATA(87)",
	OutTemp       => MIMCWRITEDATA_OUT(87),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(87),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(87), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(88),
	GlitchData    => MIMCWRITEDATA88_GlitchData,
	OutSignalName => "MIMCWRITEDATA(88)",
	OutTemp       => MIMCWRITEDATA_OUT(88),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(88),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(88), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(89),
	GlitchData    => MIMCWRITEDATA89_GlitchData,
	OutSignalName => "MIMCWRITEDATA(89)",
	OutTemp       => MIMCWRITEDATA_OUT(89),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(89),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(89), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(90),
	GlitchData    => MIMCWRITEDATA90_GlitchData,
	OutSignalName => "MIMCWRITEDATA(90)",
	OutTemp       => MIMCWRITEDATA_OUT(90),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(90),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(90), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(91),
	GlitchData    => MIMCWRITEDATA91_GlitchData,
	OutSignalName => "MIMCWRITEDATA(91)",
	OutTemp       => MIMCWRITEDATA_OUT(91),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(91),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(91), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(92),
	GlitchData    => MIMCWRITEDATA92_GlitchData,
	OutSignalName => "MIMCWRITEDATA(92)",
	OutTemp       => MIMCWRITEDATA_OUT(92),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(92),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(92), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(93),
	GlitchData    => MIMCWRITEDATA93_GlitchData,
	OutSignalName => "MIMCWRITEDATA(93)",
	OutTemp       => MIMCWRITEDATA_OUT(93),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(93),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(93), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(94),
	GlitchData    => MIMCWRITEDATA94_GlitchData,
	OutSignalName => "MIMCWRITEDATA(94)",
	OutTemp       => MIMCWRITEDATA_OUT(94),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(94),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(94), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(95),
	GlitchData    => MIMCWRITEDATA95_GlitchData,
	OutSignalName => "MIMCWRITEDATA(95)",
	OutTemp       => MIMCWRITEDATA_OUT(95),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(95),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(95), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(96),
	GlitchData    => MIMCWRITEDATA96_GlitchData,
	OutSignalName => "MIMCWRITEDATA(96)",
	OutTemp       => MIMCWRITEDATA_OUT(96),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(96),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(96), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(97),
	GlitchData    => MIMCWRITEDATA97_GlitchData,
	OutSignalName => "MIMCWRITEDATA(97)",
	OutTemp       => MIMCWRITEDATA_OUT(97),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(97),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(97), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(98),
	GlitchData    => MIMCWRITEDATA98_GlitchData,
	OutSignalName => "MIMCWRITEDATA(98)",
	OutTemp       => MIMCWRITEDATA_OUT(98),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(98),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(98), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(99),
	GlitchData    => MIMCWRITEDATA99_GlitchData,
	OutSignalName => "MIMCWRITEDATA(99)",
	OutTemp       => MIMCWRITEDATA_OUT(99),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(99),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(99), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(100),
	GlitchData    => MIMCWRITEDATA100_GlitchData,
	OutSignalName => "MIMCWRITEDATA(100)",
	OutTemp       => MIMCWRITEDATA_OUT(100),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(100),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(100), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(101),
	GlitchData    => MIMCWRITEDATA101_GlitchData,
	OutSignalName => "MIMCWRITEDATA(101)",
	OutTemp       => MIMCWRITEDATA_OUT(101),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(101),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(101), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(102),
	GlitchData    => MIMCWRITEDATA102_GlitchData,
	OutSignalName => "MIMCWRITEDATA(102)",
	OutTemp       => MIMCWRITEDATA_OUT(102),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(102),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(102), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(103),
	GlitchData    => MIMCWRITEDATA103_GlitchData,
	OutSignalName => "MIMCWRITEDATA(103)",
	OutTemp       => MIMCWRITEDATA_OUT(103),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(103),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(103), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(104),
	GlitchData    => MIMCWRITEDATA104_GlitchData,
	OutSignalName => "MIMCWRITEDATA(104)",
	OutTemp       => MIMCWRITEDATA_OUT(104),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(104),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(104), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(105),
	GlitchData    => MIMCWRITEDATA105_GlitchData,
	OutSignalName => "MIMCWRITEDATA(105)",
	OutTemp       => MIMCWRITEDATA_OUT(105),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(105),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(105), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(106),
	GlitchData    => MIMCWRITEDATA106_GlitchData,
	OutSignalName => "MIMCWRITEDATA(106)",
	OutTemp       => MIMCWRITEDATA_OUT(106),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(106),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(106), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(107),
	GlitchData    => MIMCWRITEDATA107_GlitchData,
	OutSignalName => "MIMCWRITEDATA(107)",
	OutTemp       => MIMCWRITEDATA_OUT(107),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(107),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(107), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(108),
	GlitchData    => MIMCWRITEDATA108_GlitchData,
	OutSignalName => "MIMCWRITEDATA(108)",
	OutTemp       => MIMCWRITEDATA_OUT(108),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(108),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(108), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(109),
	GlitchData    => MIMCWRITEDATA109_GlitchData,
	OutSignalName => "MIMCWRITEDATA(109)",
	OutTemp       => MIMCWRITEDATA_OUT(109),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(109),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(109), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(110),
	GlitchData    => MIMCWRITEDATA110_GlitchData,
	OutSignalName => "MIMCWRITEDATA(110)",
	OutTemp       => MIMCWRITEDATA_OUT(110),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(110),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(110), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(111),
	GlitchData    => MIMCWRITEDATA111_GlitchData,
	OutSignalName => "MIMCWRITEDATA(111)",
	OutTemp       => MIMCWRITEDATA_OUT(111),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(111),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(111), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(112),
	GlitchData    => MIMCWRITEDATA112_GlitchData,
	OutSignalName => "MIMCWRITEDATA(112)",
	OutTemp       => MIMCWRITEDATA_OUT(112),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(112),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(112), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(113),
	GlitchData    => MIMCWRITEDATA113_GlitchData,
	OutSignalName => "MIMCWRITEDATA(113)",
	OutTemp       => MIMCWRITEDATA_OUT(113),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(113),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(113), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(114),
	GlitchData    => MIMCWRITEDATA114_GlitchData,
	OutSignalName => "MIMCWRITEDATA(114)",
	OutTemp       => MIMCWRITEDATA_OUT(114),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(114),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(114), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(115),
	GlitchData    => MIMCWRITEDATA115_GlitchData,
	OutSignalName => "MIMCWRITEDATA(115)",
	OutTemp       => MIMCWRITEDATA_OUT(115),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(115),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(115), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(116),
	GlitchData    => MIMCWRITEDATA116_GlitchData,
	OutSignalName => "MIMCWRITEDATA(116)",
	OutTemp       => MIMCWRITEDATA_OUT(116),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(116),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(116), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(117),
	GlitchData    => MIMCWRITEDATA117_GlitchData,
	OutSignalName => "MIMCWRITEDATA(117)",
	OutTemp       => MIMCWRITEDATA_OUT(117),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(117),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(117), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(118),
	GlitchData    => MIMCWRITEDATA118_GlitchData,
	OutSignalName => "MIMCWRITEDATA(118)",
	OutTemp       => MIMCWRITEDATA_OUT(118),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(118),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(118), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(119),
	GlitchData    => MIMCWRITEDATA119_GlitchData,
	OutSignalName => "MIMCWRITEDATA(119)",
	OutTemp       => MIMCWRITEDATA_OUT(119),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(119),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(119), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(120),
	GlitchData    => MIMCWRITEDATA120_GlitchData,
	OutSignalName => "MIMCWRITEDATA(120)",
	OutTemp       => MIMCWRITEDATA_OUT(120),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(120),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(120), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(121),
	GlitchData    => MIMCWRITEDATA121_GlitchData,
	OutSignalName => "MIMCWRITEDATA(121)",
	OutTemp       => MIMCWRITEDATA_OUT(121),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(121),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(121), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(122),
	GlitchData    => MIMCWRITEDATA122_GlitchData,
	OutSignalName => "MIMCWRITEDATA(122)",
	OutTemp       => MIMCWRITEDATA_OUT(122),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(122),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(122), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(123),
	GlitchData    => MIMCWRITEDATA123_GlitchData,
	OutSignalName => "MIMCWRITEDATA(123)",
	OutTemp       => MIMCWRITEDATA_OUT(123),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(123),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(123), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(124),
	GlitchData    => MIMCWRITEDATA124_GlitchData,
	OutSignalName => "MIMCWRITEDATA(124)",
	OutTemp       => MIMCWRITEDATA_OUT(124),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(124),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(124), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(125),
	GlitchData    => MIMCWRITEDATA125_GlitchData,
	OutSignalName => "MIMCWRITEDATA(125)",
	OutTemp       => MIMCWRITEDATA_OUT(125),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(125),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(125), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(126),
	GlitchData    => MIMCWRITEDATA126_GlitchData,
	OutSignalName => "MIMCWRITEDATA(126)",
	OutTemp       => MIMCWRITEDATA_OUT(126),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(126),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(126), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATA(127),
	GlitchData    => MIMCWRITEDATA127_GlitchData,
	OutSignalName => "MIMCWRITEDATA(127)",
	OutTemp       => MIMCWRITEDATA_OUT(127),
	Paths       => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATA(127),TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATA(127), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => MIMCWRITEDATAVALID,
	GlitchData    => MIMCWRITEDATAVALID_GlitchData,
	OutSignalName => "MIMCWRITEDATAVALID",
	OutTemp       => MIMCWRITEDATAVALID_OUT,
	Paths         => (0 => (CPMMCCLK_dly'last_event, tpd_CPMMCCLK_MIMCWRITEDATAVALID,TRUE)),
	 DefaultDelay =>  tpd_CPMMCCLK_MIMCWRITEDATAVALID, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCCPMINTERCONNECTBUSY,
	GlitchData    => PPCCPMINTERCONNECTBUSY_GlitchData,
	OutSignalName => "PPCCPMINTERCONNECTBUSY",
	OutTemp       => PPCCPMINTERCONNECTBUSY_OUT,
	Paths         => (0 => (CPMINTERCONNECTCLK_dly'last_event, tpd_CPMINTERCONNECTCLK_PPCCPMINTERCONNECTBUSY,TRUE)),
	 DefaultDelay =>  tpd_CPMINTERCONNECTCLK_PPCCPMINTERCONNECTBUSY, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRACK,
	GlitchData    => PPCDSDCRACK_GlitchData,
	OutSignalName => "PPCDSDCRACK",
	OutTemp       => PPCDSDCRACK_OUT,
	Paths         => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRACK,TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRACK, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRTIMEOUTWAIT,
	GlitchData    => PPCDSDCRTIMEOUTWAIT_GlitchData,
	OutSignalName => "PPCDSDCRTIMEOUTWAIT",
	OutTemp       => PPCDSDCRTIMEOUTWAIT_OUT,
	Paths         => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRTIMEOUTWAIT,TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRTIMEOUTWAIT, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(0),
	GlitchData    => PPCDSDCRDBUSIN0_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(0)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(0),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(0),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(0), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(1),
	GlitchData    => PPCDSDCRDBUSIN1_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(1)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(1),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(1),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(1), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(2),
	GlitchData    => PPCDSDCRDBUSIN2_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(2)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(2),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(2),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(2), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(3),
	GlitchData    => PPCDSDCRDBUSIN3_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(3)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(3),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(3),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(3), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(4),
	GlitchData    => PPCDSDCRDBUSIN4_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(4)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(4),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(4),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(4), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(5),
	GlitchData    => PPCDSDCRDBUSIN5_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(5)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(5),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(5),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(5), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(6),
	GlitchData    => PPCDSDCRDBUSIN6_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(6)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(6),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(6),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(6), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(7),
	GlitchData    => PPCDSDCRDBUSIN7_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(7)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(7),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(7),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(7), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(8),
	GlitchData    => PPCDSDCRDBUSIN8_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(8)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(8),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(8),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(8), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(9),
	GlitchData    => PPCDSDCRDBUSIN9_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(9)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(9),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(9),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(9), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(10),
	GlitchData    => PPCDSDCRDBUSIN10_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(10)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(10),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(10),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(10), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(11),
	GlitchData    => PPCDSDCRDBUSIN11_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(11)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(11),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(11),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(11), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(12),
	GlitchData    => PPCDSDCRDBUSIN12_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(12)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(12),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(12),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(12), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(13),
	GlitchData    => PPCDSDCRDBUSIN13_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(13)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(13),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(13),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(13), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(14),
	GlitchData    => PPCDSDCRDBUSIN14_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(14)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(14),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(14),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(14), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(15),
	GlitchData    => PPCDSDCRDBUSIN15_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(15)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(15),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(15),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(15), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(16),
	GlitchData    => PPCDSDCRDBUSIN16_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(16)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(16),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(16),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(16), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(17),
	GlitchData    => PPCDSDCRDBUSIN17_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(17)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(17),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(17),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(17), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(18),
	GlitchData    => PPCDSDCRDBUSIN18_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(18)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(18),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(18),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(18), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(19),
	GlitchData    => PPCDSDCRDBUSIN19_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(19)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(19),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(19),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(19), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(20),
	GlitchData    => PPCDSDCRDBUSIN20_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(20)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(20),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(20),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(20), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(21),
	GlitchData    => PPCDSDCRDBUSIN21_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(21)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(21),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(21),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(21), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(22),
	GlitchData    => PPCDSDCRDBUSIN22_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(22)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(22),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(22),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(22), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(23),
	GlitchData    => PPCDSDCRDBUSIN23_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(23)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(23),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(23),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(23), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(24),
	GlitchData    => PPCDSDCRDBUSIN24_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(24)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(24),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(24),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(24), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(25),
	GlitchData    => PPCDSDCRDBUSIN25_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(25)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(25),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(25),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(25), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(26),
	GlitchData    => PPCDSDCRDBUSIN26_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(26)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(26),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(26),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(26), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(27),
	GlitchData    => PPCDSDCRDBUSIN27_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(27)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(27),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(27),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(27), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(28),
	GlitchData    => PPCDSDCRDBUSIN28_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(28)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(28),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(28),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(28), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(29),
	GlitchData    => PPCDSDCRDBUSIN29_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(29)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(29),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(29),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(29), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(30),
	GlitchData    => PPCDSDCRDBUSIN30_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(30)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(30),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(30),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(30), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCDSDCRDBUSIN(31),
	GlitchData    => PPCDSDCRDBUSIN31_GlitchData,
	OutSignalName => "PPCDSDCRDBUSIN(31)",
	OutTemp       => PPCDSDCRDBUSIN_OUT(31),
	Paths       => (0 => (CPMDCRCLK_dly'last_event, tpd_CPMDCRCLK_PPCDSDCRDBUSIN(31),TRUE)),
	 DefaultDelay =>  tpd_CPMDCRCLK_PPCDSDCRDBUSIN(31), 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);
	VitalPathDelay01
	(
	OutSignal     => PPCEICINTERCONNECTIRQ,
	GlitchData    => PPCEICINTERCONNECTIRQ_GlitchData,
	OutSignalName => "PPCEICINTERCONNECTIRQ",
	OutTemp       => PPCEICINTERCONNECTIRQ_OUT,
	Paths         => (0 => (CPMINTERCONNECTCLK_dly'last_event, tpd_CPMINTERCONNECTCLK_PPCEICINTERCONNECTIRQ,TRUE)),
	 DefaultDelay =>  tpd_CPMINTERCONNECTCLK_PPCEICINTERCONNECTIRQ, 
	Mode          => VitalTransport,
	Xon           => false,
	MsgOn         => false,
	MsgSeverity   => WARNING
	);

   wait on
	APUFCMDECFPUOP_out,
	APUFCMDECLDSTXFERSIZE_out,
	APUFCMDECLOAD_out,
	APUFCMDECNONAUTON_out,
	APUFCMDECSTORE_out,
	APUFCMDECUDIVALID_out,
	APUFCMDECUDI_out,
	APUFCMENDIAN_out,
	APUFCMFLUSH_out,
	APUFCMINSTRUCTION_out,
	APUFCMINSTRVALID_out,
	APUFCMLOADBYTEADDR_out,
	APUFCMLOADDATA_out,
	APUFCMLOADDVALID_out,
	APUFCMMSRFE0_out,
	APUFCMMSRFE1_out,
	APUFCMNEXTINSTRREADY_out,
	APUFCMOPERANDVALID_out,
	APUFCMRADATA_out,
	APUFCMRBDATA_out,
	APUFCMWRITEBACKOK_out,
	C440CPMCORESLEEPREQ_out,
	C440CPMDECIRPTREQ_out,
	C440CPMFITIRPTREQ_out,
	C440CPMMSRCE_out,
	C440CPMMSREE_out,
	C440CPMTIMERRESETREQ_out,
	C440CPMWDIRPTREQ_out,
	C440DBGSYSTEMCONTROL_out,
	C440JTGTDOEN_out,
	C440JTGTDO_out,
	C440MACHINECHECK_out,
	C440RSTCHIPRESETREQ_out,
	C440RSTCORERESETREQ_out,
	C440RSTSYSTEMRESETREQ_out,
	C440TRCBRANCHSTATUS_out,
	C440TRCCYCLE_out,
	C440TRCEXECUTIONSTATUS_out,
	C440TRCTRACESTATUS_out,
	C440TRCTRIGGEREVENTOUT_out,
	C440TRCTRIGGEREVENTTYPE_out,
	DMA0LLRSTENGINEACK_out,
	DMA0LLRXDSTRDYN_out,
	DMA0LLTXD_out,
	DMA0LLTXEOFN_out,
	DMA0LLTXEOPN_out,
	DMA0LLTXREM_out,
	DMA0LLTXSOFN_out,
	DMA0LLTXSOPN_out,
	DMA0LLTXSRCRDYN_out,
	DMA0RXIRQ_out,
	DMA0TXIRQ_out,
	DMA1LLRSTENGINEACK_out,
	DMA1LLRXDSTRDYN_out,
	DMA1LLTXD_out,
	DMA1LLTXEOFN_out,
	DMA1LLTXEOPN_out,
	DMA1LLTXREM_out,
	DMA1LLTXSOFN_out,
	DMA1LLTXSOPN_out,
	DMA1LLTXSRCRDYN_out,
	DMA1RXIRQ_out,
	DMA1TXIRQ_out,
	DMA2LLRSTENGINEACK_out,
	DMA2LLRXDSTRDYN_out,
	DMA2LLTXD_out,
	DMA2LLTXEOFN_out,
	DMA2LLTXEOPN_out,
	DMA2LLTXREM_out,
	DMA2LLTXSOFN_out,
	DMA2LLTXSOPN_out,
	DMA2LLTXSRCRDYN_out,
	DMA2RXIRQ_out,
	DMA2TXIRQ_out,
	DMA3LLRSTENGINEACK_out,
	DMA3LLRXDSTRDYN_out,
	DMA3LLTXD_out,
	DMA3LLTXEOFN_out,
	DMA3LLTXEOPN_out,
	DMA3LLTXREM_out,
	DMA3LLTXSOFN_out,
	DMA3LLTXSOPN_out,
	DMA3LLTXSRCRDYN_out,
	DMA3RXIRQ_out,
	DMA3TXIRQ_out,
	MIMCADDRESSVALID_out,
	MIMCADDRESS_out,
	MIMCBANKCONFLICT_out,
	MIMCBYTEENABLE_out,
	MIMCREADNOTWRITE_out,
	MIMCROWCONFLICT_out,
	MIMCWRITEDATAVALID_out,
	MIMCWRITEDATA_out,
	PPCCPMINTERCONNECTBUSY_out,
	PPCDMDCRABUS_out,
	PPCDMDCRDBUSOUT_out,
	PPCDMDCRREAD_out,
	PPCDMDCRUABUS_out,
	PPCDMDCRWRITE_out,
	PPCDSDCRACK_out,
	PPCDSDCRDBUSIN_out,
	PPCDSDCRTIMEOUTWAIT_out,
	PPCEICINTERCONNECTIRQ_out,
	PPCMPLBABORT_out,
	PPCMPLBABUS_out,
	PPCMPLBBE_out,
	PPCMPLBBUSLOCK_out,
	PPCMPLBLOCKERR_out,
	PPCMPLBPRIORITY_out,
	PPCMPLBRDBURST_out,
	PPCMPLBREQUEST_out,
	PPCMPLBRNW_out,
	PPCMPLBSIZE_out,
	PPCMPLBTATTRIBUTE_out,
	PPCMPLBTYPE_out,
	PPCMPLBUABUS_out,
	PPCMPLBWRBURST_out,
	PPCMPLBWRDBUS_out,
	PPCS0PLBADDRACK_out,
	PPCS0PLBMBUSY_out,
	PPCS0PLBMIRQ_out,
	PPCS0PLBMRDERR_out,
	PPCS0PLBMWRERR_out,
	PPCS0PLBRDBTERM_out,
	PPCS0PLBRDCOMP_out,
	PPCS0PLBRDDACK_out,
	PPCS0PLBRDDBUS_out,
	PPCS0PLBRDWDADDR_out,
	PPCS0PLBREARBITRATE_out,
	PPCS0PLBSSIZE_out,
	PPCS0PLBWAIT_out,
	PPCS0PLBWRBTERM_out,
	PPCS0PLBWRCOMP_out,
	PPCS0PLBWRDACK_out,
	PPCS1PLBADDRACK_out,
	PPCS1PLBMBUSY_out,
	PPCS1PLBMIRQ_out,
	PPCS1PLBMRDERR_out,
	PPCS1PLBMWRERR_out,
	PPCS1PLBRDBTERM_out,
	PPCS1PLBRDCOMP_out,
	PPCS1PLBRDDACK_out,
	PPCS1PLBRDDBUS_out,
	PPCS1PLBRDWDADDR_out,
	PPCS1PLBREARBITRATE_out,
	PPCS1PLBSSIZE_out,
	PPCS1PLBWAIT_out,
	PPCS1PLBWRBTERM_out,
	PPCS1PLBWRCOMP_out,
	PPCS1PLBWRDACK_out,

	CPMC440CORECLOCKINACTIVE_dly,
	CPMINTERCONNECTCLKNTO1_dly,
	DBGC440DEBUGHALT_dly,
	DBGC440SYSTEMSTATUS_dly,
	DBGC440UNCONDDEBUGEVENT_dly,
	DCRPPCDMACK_dly,
	DCRPPCDMDBUSIN_dly,
	DCRPPCDMTIMEOUTWAIT_dly,
	DCRPPCDSABUS_dly,
	DCRPPCDSDBUSOUT_dly,
	DCRPPCDSREAD_dly,
	DCRPPCDSWRITE_dly,
	FCMAPUCONFIRMINSTR_dly,
	FCMAPUCR_dly,
	FCMAPUDONE_dly,
	FCMAPUEXCEPTION_dly,
	FCMAPUFPSCRFEX_dly,
	FCMAPURESULTVALID_dly,
	FCMAPURESULT_dly,
	FCMAPUSLEEPNOTREADY_dly,
	FCMAPUSTOREDATA_dly,
	JTGC440TDI_dly,
	JTGC440TMS_dly,
	LLDMA0RSTENGINEREQ_dly,
	LLDMA0RXD_dly,
	LLDMA0RXEOFN_dly,
	LLDMA0RXEOPN_dly,
	LLDMA0RXREM_dly,
	LLDMA0RXSOFN_dly,
	LLDMA0RXSOPN_dly,
	LLDMA0RXSRCRDYN_dly,
	LLDMA0TXDSTRDYN_dly,
	LLDMA1RSTENGINEREQ_dly,
	LLDMA1RXD_dly,
	LLDMA1RXEOFN_dly,
	LLDMA1RXEOPN_dly,
	LLDMA1RXREM_dly,
	LLDMA1RXSOFN_dly,
	LLDMA1RXSOPN_dly,
	LLDMA1RXSRCRDYN_dly,
	LLDMA1TXDSTRDYN_dly,
	LLDMA2RSTENGINEREQ_dly,
	LLDMA2RXD_dly,
	LLDMA2RXEOFN_dly,
	LLDMA2RXEOPN_dly,
	LLDMA2RXREM_dly,
	LLDMA2RXSOFN_dly,
	LLDMA2RXSOPN_dly,
	LLDMA2RXSRCRDYN_dly,
	LLDMA2TXDSTRDYN_dly,
	LLDMA3RSTENGINEREQ_dly,
	LLDMA3RXD_dly,
	LLDMA3RXEOFN_dly,
	LLDMA3RXEOPN_dly,
	LLDMA3RXREM_dly,
	LLDMA3RXSOFN_dly,
	LLDMA3RXSOPN_dly,
	LLDMA3RXSRCRDYN_dly,
	LLDMA3TXDSTRDYN_dly,
	MCMIADDRREADYTOACCEPT_dly,
	MCMIREADDATAERR_dly,
	MCMIREADDATAVALID_dly,
	MCMIREADDATA_dly,
	PLBPPCMADDRACK_dly,
	PLBPPCMMBUSY_dly,
	PLBPPCMMIRQ_dly,
	PLBPPCMMRDERR_dly,
	PLBPPCMMWRERR_dly,
	PLBPPCMRDBTERM_dly,
	PLBPPCMRDDACK_dly,
	PLBPPCMRDDBUS_dly,
	PLBPPCMRDPENDPRI_dly,
	PLBPPCMRDPENDREQ_dly,
	PLBPPCMRDWDADDR_dly,
	PLBPPCMREARBITRATE_dly,
	PLBPPCMREQPRI_dly,
	PLBPPCMSSIZE_dly,
	PLBPPCMTIMEOUT_dly,
	PLBPPCMWRBTERM_dly,
	PLBPPCMWRDACK_dly,
	PLBPPCMWRPENDPRI_dly,
	PLBPPCMWRPENDREQ_dly,
	PLBPPCS0ABORT_dly,
	PLBPPCS0ABUS_dly,
	PLBPPCS0BE_dly,
	PLBPPCS0BUSLOCK_dly,
	PLBPPCS0LOCKERR_dly,
	PLBPPCS0MASTERID_dly,
	PLBPPCS0MSIZE_dly,
	PLBPPCS0PAVALID_dly,
	PLBPPCS0RDBURST_dly,
	PLBPPCS0RDPENDPRI_dly,
	PLBPPCS0RDPENDREQ_dly,
	PLBPPCS0RDPRIM_dly,
	PLBPPCS0REQPRI_dly,
	PLBPPCS0RNW_dly,
	PLBPPCS0SAVALID_dly,
	PLBPPCS0SIZE_dly,
	PLBPPCS0TATTRIBUTE_dly,
	PLBPPCS0TYPE_dly,
	PLBPPCS0UABUS_dly,
	PLBPPCS0WRBURST_dly,
	PLBPPCS0WRDBUS_dly,
	PLBPPCS0WRPENDPRI_dly,
	PLBPPCS0WRPENDREQ_dly,
	PLBPPCS0WRPRIM_dly,
	PLBPPCS1ABORT_dly,
	PLBPPCS1ABUS_dly,
	PLBPPCS1BE_dly,
	PLBPPCS1BUSLOCK_dly,
	PLBPPCS1LOCKERR_dly,
	PLBPPCS1MASTERID_dly,
	PLBPPCS1MSIZE_dly,
	PLBPPCS1PAVALID_dly,
	PLBPPCS1RDBURST_dly,
	PLBPPCS1RDPENDPRI_dly,
	PLBPPCS1RDPENDREQ_dly,
	PLBPPCS1RDPRIM_dly,
	PLBPPCS1REQPRI_dly,
	PLBPPCS1RNW_dly,
	PLBPPCS1SAVALID_dly,
	PLBPPCS1SIZE_dly,
	PLBPPCS1TATTRIBUTE_dly,
	PLBPPCS1TYPE_dly,
	PLBPPCS1UABUS_dly,
	PLBPPCS1WRBURST_dly,
	PLBPPCS1WRDBUS_dly,
	PLBPPCS1WRPENDPRI_dly,
	PLBPPCS1WRPENDREQ_dly,
	PLBPPCS1WRPRIM_dly,
	TRCC440TRACEDISABLE_dly,
	TRCC440TRIGGEREVENTIN_dly;

	end process TIMING;

end X_PPC440_V;
